
module DADDA_16x16_42 ( a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [31:0] out;
  wire   add_168_CI, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1118, n1120, n1122, n1124, n1126, n1128, n1130,
         n1132, n1134, n1136, n1138, n1140, n1142, n1144, n1146, n1148, n1149,
         n1151, n1153, n1155, n1157, n1159, n1161, n1163, n1165, n1167, n1169,
         n1171, n1173, n1174, n1176, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237;
  wire   [255:1] p;
  wire   [111:84] s;
  wire   [110:84] c;

  FAxp33_ASAP7_6t_L add_168_U1_0 ( .A(p[1]), .B(p[16]), .CI(add_168_CI), .CON(
        n1179), .SN(n1178) );
  FAxp33_ASAP7_6t_L add_168_U1_1 ( .A(s[84]), .B(p[32]), .CI(n1176), .CON(
        n1181), .SN(n1180) );
  FAxp33_ASAP7_6t_L add_168_U1_2 ( .A(n1173), .B(c[84]), .CI(n1174), .CON(
        n1183), .SN(n1182) );
  FAxp33_ASAP7_6t_L add_168_U1_3 ( .A(s[86]), .B(c[85]), .CI(n1171), .CON(
        n1185), .SN(n1184) );
  FAxp33_ASAP7_6t_L add_168_U1_4 ( .A(s[87]), .B(c[86]), .CI(n1169), .CON(
        n1187), .SN(n1186) );
  FAxp33_ASAP7_6t_L add_168_U1_5 ( .A(s[88]), .B(c[87]), .CI(n1167), .CON(
        n1189), .SN(n1188) );
  FAxp33_ASAP7_6t_L add_168_U1_6 ( .A(s[89]), .B(c[88]), .CI(n1165), .CON(
        n1191), .SN(n1190) );
  FAxp33_ASAP7_6t_L add_168_U1_7 ( .A(s[90]), .B(c[89]), .CI(n1163), .CON(
        n1193), .SN(n1192) );
  FAxp33_ASAP7_6t_L add_168_U1_8 ( .A(s[91]), .B(c[90]), .CI(n1161), .CON(
        n1195), .SN(n1194) );
  FAxp33_ASAP7_6t_L add_168_U1_9 ( .A(s[92]), .B(c[91]), .CI(n1159), .CON(
        n1197), .SN(n1196) );
  FAxp33_ASAP7_6t_L add_168_U1_10 ( .A(s[93]), .B(c[92]), .CI(n1157), .CON(
        n1199), .SN(n1198) );
  FAxp33_ASAP7_6t_L add_168_U1_11 ( .A(s[94]), .B(c[93]), .CI(n1155), .CON(
        n1201), .SN(n1200) );
  FAxp33_ASAP7_6t_L add_168_U1_12 ( .A(s[95]), .B(c[94]), .CI(n1153), .CON(
        n1203), .SN(n1202) );
  FAxp33_ASAP7_6t_L add_168_U1_13 ( .A(s[96]), .B(c[95]), .CI(n1151), .CON(
        n1205), .SN(n1204) );
  FAxp33_ASAP7_6t_L add_168_U1_14 ( .A(s[97]), .B(c[96]), .CI(n1149), .CON(
        n1207), .SN(n1206) );
  FAxp33_ASAP7_6t_L add_168_U1_15 ( .A(s[98]), .B(c[97]), .CI(n1146), .CON(
        n1209), .SN(n1208) );
  FAxp33_ASAP7_6t_L add_168_U1_16 ( .A(s[99]), .B(c[98]), .CI(n1144), .CON(
        n1211), .SN(n1210) );
  FAxp33_ASAP7_6t_L add_168_U1_17 ( .A(s[100]), .B(c[99]), .CI(n1142), .CON(
        n1213), .SN(n1212) );
  FAxp33_ASAP7_6t_L add_168_U1_18 ( .A(s[101]), .B(c[100]), .CI(n1140), .CON(
        n1215), .SN(n1214) );
  FAxp33_ASAP7_6t_L add_168_U1_19 ( .A(s[102]), .B(c[101]), .CI(n1138), .CON(
        n1217), .SN(n1216) );
  FAxp33_ASAP7_6t_L add_168_U1_20 ( .A(s[103]), .B(c[102]), .CI(n1136), .CON(
        n1219), .SN(n1218) );
  FAxp33_ASAP7_6t_L add_168_U1_21 ( .A(s[104]), .B(c[103]), .CI(n1134), .CON(
        n1221), .SN(n1220) );
  FAxp33_ASAP7_6t_L add_168_U1_22 ( .A(s[105]), .B(c[104]), .CI(n1132), .CON(
        n1223), .SN(n1222) );
  FAxp33_ASAP7_6t_L add_168_U1_23 ( .A(s[106]), .B(c[105]), .CI(n1130), .CON(
        n1225), .SN(n1224) );
  FAxp33_ASAP7_6t_L add_168_U1_24 ( .A(s[107]), .B(c[106]), .CI(n1128), .CON(
        n1227), .SN(n1226) );
  FAxp33_ASAP7_6t_L add_168_U1_25 ( .A(s[108]), .B(c[107]), .CI(n1126), .CON(
        n1229), .SN(n1228) );
  FAxp33_ASAP7_6t_L add_168_U1_26 ( .A(s[109]), .B(c[108]), .CI(n1124), .CON(
        n1231), .SN(n1230) );
  FAxp33_ASAP7_6t_L add_168_U1_27 ( .A(s[110]), .B(c[109]), .CI(n1122), .CON(
        n1233), .SN(n1232) );
  FAxp33_ASAP7_6t_L add_168_U1_28 ( .A(s[111]), .B(c[110]), .CI(n1120), .CON(
        n1235), .SN(n1234) );
  FAxp33_ASAP7_6t_L add_168_U1_29 ( .A(p[255]), .B(n1148), .CI(n1118), .CON(
        n1237), .SN(n1236) );
  TIELOxp5_ASAP7_6t_L U292 ( .L(add_168_CI) );
  XOR2xp5r_ASAP7_6t_L U293 ( .A(n35), .B(n36), .Y(s[99]) );
  XOR2xp5r_ASAP7_6t_L U294 ( .A(n37), .B(n38), .Y(s[98]) );
  XOR2xp5r_ASAP7_6t_L U295 ( .A(n39), .B(n40), .Y(s[97]) );
  XOR2xp5r_ASAP7_6t_L U296 ( .A(n41), .B(n42), .Y(s[96]) );
  XOR2xp5r_ASAP7_6t_L U297 ( .A(n43), .B(n44), .Y(s[95]) );
  XOR2xp5r_ASAP7_6t_L U298 ( .A(n45), .B(n46), .Y(s[94]) );
  XOR2xp5r_ASAP7_6t_L U299 ( .A(n47), .B(n48), .Y(s[93]) );
  XOR2xp5r_ASAP7_6t_L U300 ( .A(n49), .B(n50), .Y(s[92]) );
  XOR2xp5r_ASAP7_6t_L U301 ( .A(n51), .B(n52), .Y(s[91]) );
  XOR2xp5r_ASAP7_6t_L U302 ( .A(n53), .B(n54), .Y(s[90]) );
  XOR2xp5r_ASAP7_6t_L U303 ( .A(n55), .B(n56), .Y(s[89]) );
  XOR2xp5r_ASAP7_6t_L U304 ( .A(n57), .B(n58), .Y(s[88]) );
  XOR2xp5r_ASAP7_6t_L U305 ( .A(n59), .B(n60), .Y(s[87]) );
  XOR2xp5r_ASAP7_6t_L U306 ( .A(n61), .B(n62), .Y(s[86]) );
  XOR2xp5r_ASAP7_6t_L U307 ( .A(n63), .B(n64), .Y(s[84]) );
  NAND2xp5R_ASAP7_6t_L U308 ( .A(a[1]), .B(b[1]), .Y(n63) );
  XOR2xp5r_ASAP7_6t_L U309 ( .A(n65), .B(n66), .Y(s[111]) );
  XOR2xp5r_ASAP7_6t_L U310 ( .A(n67), .B(n68), .Y(s[110]) );
  XOR2xp5r_ASAP7_6t_L U311 ( .A(n69), .B(n70), .Y(s[109]) );
  XOR2xp5r_ASAP7_6t_L U312 ( .A(n71), .B(n72), .Y(s[108]) );
  XOR2xp5r_ASAP7_6t_L U313 ( .A(n73), .B(n74), .Y(s[107]) );
  XOR2xp5r_ASAP7_6t_L U314 ( .A(n75), .B(n76), .Y(s[106]) );
  XOR2xp5r_ASAP7_6t_L U315 ( .A(n77), .B(n78), .Y(s[105]) );
  XOR2xp5r_ASAP7_6t_L U316 ( .A(n79), .B(n80), .Y(s[104]) );
  XOR2xp5r_ASAP7_6t_L U317 ( .A(n81), .B(n82), .Y(s[103]) );
  XOR2xp5r_ASAP7_6t_L U318 ( .A(n83), .B(n84), .Y(s[102]) );
  XOR2xp5r_ASAP7_6t_L U319 ( .A(n85), .B(n86), .Y(s[101]) );
  XOR2xp5r_ASAP7_6t_L U320 ( .A(n87), .B(n88), .Y(s[100]) );
  NOR2xp5_ASAP7_6t_L U321 ( .A(n89), .B(n90), .Y(p[32]) );
  NOR2xp5_ASAP7_6t_L U322 ( .A(n91), .B(n92), .Y(p[255]) );
  NOR2xp5_ASAP7_6t_L U323 ( .A(n93), .B(n94), .Y(p[1]) );
  NOR2xp5_ASAP7_6t_L U324 ( .A(n89), .B(n95), .Y(p[16]) );
  NOR2xp5_ASAP7_6t_L U325 ( .A(n89), .B(n94), .Y(out[0]) );
  INVx1_ASAP7_6t_L U326 ( .A(n1237), .Y(out[31]) );
  INVx1_ASAP7_6t_L U327 ( .A(n1236), .Y(out[30]) );
  INVx1_ASAP7_6t_L U328 ( .A(n1235), .Y(n1118) );
  INVx1_ASAP7_6t_L U329 ( .A(n1234), .Y(out[29]) );
  INVx1_ASAP7_6t_L U330 ( .A(n1233), .Y(n1120) );
  INVx1_ASAP7_6t_L U331 ( .A(n1232), .Y(out[28]) );
  INVx1_ASAP7_6t_L U332 ( .A(n1231), .Y(n1122) );
  INVx1_ASAP7_6t_L U333 ( .A(n1230), .Y(out[27]) );
  INVx1_ASAP7_6t_L U334 ( .A(n1229), .Y(n1124) );
  INVx1_ASAP7_6t_L U335 ( .A(n1228), .Y(out[26]) );
  INVx1_ASAP7_6t_L U336 ( .A(n1227), .Y(n1126) );
  INVx1_ASAP7_6t_L U337 ( .A(n1226), .Y(out[25]) );
  INVx1_ASAP7_6t_L U338 ( .A(n1225), .Y(n1128) );
  INVx1_ASAP7_6t_L U339 ( .A(n1224), .Y(out[24]) );
  INVx1_ASAP7_6t_L U340 ( .A(n1223), .Y(n1130) );
  INVx1_ASAP7_6t_L U341 ( .A(n1222), .Y(out[23]) );
  INVx1_ASAP7_6t_L U342 ( .A(n1221), .Y(n1132) );
  INVx1_ASAP7_6t_L U343 ( .A(n1220), .Y(out[22]) );
  INVx1_ASAP7_6t_L U344 ( .A(n1219), .Y(n1134) );
  INVx1_ASAP7_6t_L U345 ( .A(n1218), .Y(out[21]) );
  INVx1_ASAP7_6t_L U346 ( .A(n1217), .Y(n1136) );
  INVx1_ASAP7_6t_L U347 ( .A(n1216), .Y(out[20]) );
  INVx1_ASAP7_6t_L U348 ( .A(n1215), .Y(n1138) );
  INVx1_ASAP7_6t_L U349 ( .A(n1214), .Y(out[19]) );
  INVx1_ASAP7_6t_L U350 ( .A(n1213), .Y(n1140) );
  INVx1_ASAP7_6t_L U351 ( .A(n1212), .Y(out[18]) );
  INVx1_ASAP7_6t_L U352 ( .A(n1211), .Y(n1142) );
  INVx1_ASAP7_6t_L U353 ( .A(n1210), .Y(out[17]) );
  INVx1_ASAP7_6t_L U354 ( .A(n1209), .Y(n1144) );
  INVx1_ASAP7_6t_L U355 ( .A(n1208), .Y(out[16]) );
  INVx1_ASAP7_6t_L U356 ( .A(n1207), .Y(n1146) );
  INVx1_ASAP7_6t_L U357 ( .A(n1206), .Y(out[15]) );
  AO21x1_ASAP7_6t_L U358 ( .A1(n66), .A2(n65), .B(n96), .Y(n1148) );
  NOR3x1f_ASAP7_6t_L U359 ( .A(n97), .B(n91), .C(n98), .Y(n96) );
  OR2x2_ASAP7_6t_L U360 ( .A(n99), .B(n100), .Y(n65) );
  NOR3x1f_ASAP7_6t_L U361 ( .A(n101), .B(n102), .C(n92), .Y(n100) );
  NOR3x1f_ASAP7_6t_L U362 ( .A(n103), .B(n104), .C(n98), .Y(n99) );
  XOR2xp5r_ASAP7_6t_L U363 ( .A(n105), .B(n97), .Y(n66) );
  NAND2xp5R_ASAP7_6t_L U364 ( .A(b[15]), .B(a[14]), .Y(n97) );
  NAND2xp5R_ASAP7_6t_L U365 ( .A(a[15]), .B(b[14]), .Y(n105) );
  INVx1_ASAP7_6t_L U366 ( .A(n1205), .Y(n1149) );
  INVx1_ASAP7_6t_L U367 ( .A(n1204), .Y(out[14]) );
  INVx1_ASAP7_6t_L U368 ( .A(n1203), .Y(n1151) );
  INVx1_ASAP7_6t_L U369 ( .A(n1202), .Y(out[13]) );
  INVx1_ASAP7_6t_L U370 ( .A(n1201), .Y(n1153) );
  INVx1_ASAP7_6t_L U371 ( .A(n1200), .Y(out[12]) );
  INVx1_ASAP7_6t_L U372 ( .A(n1199), .Y(n1155) );
  INVx1_ASAP7_6t_L U373 ( .A(n1198), .Y(out[11]) );
  INVx1_ASAP7_6t_L U374 ( .A(n1197), .Y(n1157) );
  INVx1_ASAP7_6t_L U375 ( .A(n1196), .Y(out[10]) );
  INVx1_ASAP7_6t_L U376 ( .A(n1195), .Y(n1159) );
  INVx1_ASAP7_6t_L U377 ( .A(n1194), .Y(out[9]) );
  INVx1_ASAP7_6t_L U378 ( .A(n1193), .Y(n1161) );
  INVx1_ASAP7_6t_L U379 ( .A(n1192), .Y(out[8]) );
  INVx1_ASAP7_6t_L U380 ( .A(n1191), .Y(n1163) );
  INVx1_ASAP7_6t_L U381 ( .A(n1190), .Y(out[7]) );
  INVx1_ASAP7_6t_L U382 ( .A(n1189), .Y(n1165) );
  INVx1_ASAP7_6t_L U383 ( .A(n1188), .Y(out[6]) );
  INVx1_ASAP7_6t_L U384 ( .A(n1187), .Y(n1167) );
  INVx1_ASAP7_6t_L U385 ( .A(n1186), .Y(out[5]) );
  INVx1_ASAP7_6t_L U386 ( .A(n1185), .Y(n1169) );
  INVx1_ASAP7_6t_L U387 ( .A(n1184), .Y(out[4]) );
  INVx1_ASAP7_6t_L U388 ( .A(n1183), .Y(n1171) );
  INVx1_ASAP7_6t_L U389 ( .A(n1182), .Y(out[3]) );
  INVx1_ASAP7_6t_L U390 ( .A(n1181), .Y(n1174) );
  INVx1_ASAP7_6t_L U391 ( .A(n1180), .Y(out[2]) );
  INVx1_ASAP7_6t_L U392 ( .A(n1179), .Y(n1176) );
  INVx1_ASAP7_6t_L U393 ( .A(n1178), .Y(out[1]) );
  OAI22xp5_ASAP7_6t_L U394 ( .A1(n106), .A2(n107), .B1(n36), .B2(n35), .Y(
        c[99]) );
  AOI22xp25_ASAP7_6t_L U395 ( .A1(n108), .A2(n109), .B1(n110), .B2(n111), .Y(
        n35) );
  INVx1_ASAP7_6t_L U396 ( .A(n112), .Y(n111) );
  INVx1_ASAP7_6t_L U397 ( .A(n108), .Y(n110) );
  INVx1_ASAP7_6t_L U398 ( .A(n107), .Y(n36) );
  XOR2xp5r_ASAP7_6t_L U399 ( .A(n113), .B(n114), .Y(n107) );
  XOR2xp5r_ASAP7_6t_L U400 ( .A(n106), .B(n115), .Y(n113) );
  AOI22xp25_ASAP7_6t_L U401 ( .A1(n116), .A2(n117), .B1(n118), .B2(n119), .Y(
        n106) );
  OAI22xp5_ASAP7_6t_L U402 ( .A1(n37), .A2(n38), .B1(n120), .B2(n121), .Y(
        c[98]) );
  INVx1_ASAP7_6t_L U403 ( .A(n38), .Y(n120) );
  XOR2xp5r_ASAP7_6t_L U404 ( .A(n121), .B(n122), .Y(n38) );
  XOR2xp5r_ASAP7_6t_L U405 ( .A(n109), .B(n108), .Y(n122) );
  OAI22xp5_ASAP7_6t_L U406 ( .A1(n123), .A2(n124), .B1(n125), .B2(n126), .Y(
        n108) );
  XOR2xp5r_ASAP7_6t_L U407 ( .A(n127), .B(n112), .Y(n126) );
  XOR2xp5r_ASAP7_6t_L U408 ( .A(n128), .B(n112), .Y(n124) );
  XOR2xp5r_ASAP7_6t_L U409 ( .A(n129), .B(n130), .Y(n112) );
  XOR2xp5r_ASAP7_6t_L U410 ( .A(n116), .B(n117), .Y(n109) );
  INVx1_ASAP7_6t_L U411 ( .A(n118), .Y(n117) );
  XOR2xp5r_ASAP7_6t_L U412 ( .A(n131), .B(n132), .Y(n118) );
  XOR2xp5r_ASAP7_6t_L U413 ( .A(n119), .B(n133), .Y(n132) );
  NOR3x1f_ASAP7_6t_L U414 ( .A(n134), .B(n91), .C(n89), .Y(n119) );
  AO22x1_ASAP7_6t_L U415 ( .A1(n135), .A2(n134), .B1(n136), .B2(n137), .Y(n116) );
  INVx1_ASAP7_6t_L U416 ( .A(n136), .Y(n135) );
  AOI22xp25_ASAP7_6t_L U417 ( .A1(n138), .A2(n139), .B1(n140), .B2(n141), .Y(
        n121) );
  AOI22xp25_ASAP7_6t_L U418 ( .A1(n142), .A2(n143), .B1(n144), .B2(n145), .Y(
        n37) );
  INVx1_ASAP7_6t_L U419 ( .A(n142), .Y(n144) );
  OAI22xp5_ASAP7_6t_L U420 ( .A1(n39), .A2(n40), .B1(n146), .B2(n147), .Y(
        c[97]) );
  INVx1_ASAP7_6t_L U421 ( .A(n40), .Y(n146) );
  XOR2xp5r_ASAP7_6t_L U422 ( .A(n147), .B(n148), .Y(n40) );
  XOR2xp5r_ASAP7_6t_L U423 ( .A(n143), .B(n142), .Y(n148) );
  OAI22xp5_ASAP7_6t_L U424 ( .A1(n149), .A2(n150), .B1(n151), .B2(n152), .Y(
        n142) );
  XOR2xp5r_ASAP7_6t_L U425 ( .A(n153), .B(n145), .Y(n152) );
  XOR2xp5r_ASAP7_6t_L U426 ( .A(n154), .B(n145), .Y(n150) );
  XOR2xp5r_ASAP7_6t_L U427 ( .A(n128), .B(n125), .Y(n145) );
  INVx1_ASAP7_6t_L U428 ( .A(n123), .Y(n125) );
  XOR2xp5r_ASAP7_6t_L U429 ( .A(n155), .B(n156), .Y(n123) );
  XOR2xp5r_ASAP7_6t_L U430 ( .A(n127), .B(n157), .Y(n155) );
  OAI22xp5_ASAP7_6t_L U431 ( .A1(n158), .A2(n159), .B1(n160), .B2(n161), .Y(
        n127) );
  OAI22xp5_ASAP7_6t_L U432 ( .A1(n162), .A2(n163), .B1(n164), .B2(n165), .Y(
        n128) );
  XOR2xp5r_ASAP7_6t_L U433 ( .A(n139), .B(n138), .Y(n143) );
  AO22x1_ASAP7_6t_L U434 ( .A1(n166), .A2(n167), .B1(n168), .B2(n169), .Y(n138) );
  INVx1_ASAP7_6t_L U435 ( .A(n166), .Y(n168) );
  INVx1_ASAP7_6t_L U436 ( .A(n140), .Y(n139) );
  XOR2xp5r_ASAP7_6t_L U437 ( .A(n170), .B(n136), .Y(n140) );
  AOI22xp25_ASAP7_6t_L U438 ( .A1(n171), .A2(n172), .B1(n173), .B2(n174), .Y(
        n136) );
  XOR2xp5r_ASAP7_6t_L U439 ( .A(n175), .B(n137), .Y(n174) );
  INVx1_ASAP7_6t_L U440 ( .A(n171), .Y(n173) );
  XOR2xp5r_ASAP7_6t_L U441 ( .A(n176), .B(n137), .Y(n172) );
  XOR2xp5r_ASAP7_6t_L U442 ( .A(n177), .B(n178), .Y(n137) );
  XOR2xp5r_ASAP7_6t_L U443 ( .A(n141), .B(n134), .Y(n170) );
  XOR2xp5r_ASAP7_6t_L U444 ( .A(n179), .B(n180), .Y(n134) );
  XOR2xp5r_ASAP7_6t_L U445 ( .A(n181), .B(n182), .Y(n180) );
  NOR2xp5_ASAP7_6t_L U446 ( .A(n91), .B(n89), .Y(n181) );
  NOR3x1f_ASAP7_6t_L U447 ( .A(n183), .B(n102), .C(n93), .Y(n141) );
  AOI21xp25_ASAP7_6t_L U448 ( .A1(n184), .A2(n185), .B(n186), .Y(n147) );
  NOR3x1f_ASAP7_6t_L U449 ( .A(n184), .B(n104), .C(n89), .Y(n186) );
  AOI22xp25_ASAP7_6t_L U450 ( .A1(n187), .A2(n188), .B1(n189), .B2(n190), .Y(
        n39) );
  INVx1_ASAP7_6t_L U451 ( .A(n187), .Y(n189) );
  OAI22xp5_ASAP7_6t_L U452 ( .A1(n41), .A2(n42), .B1(n191), .B2(n192), .Y(
        c[96]) );
  INVx1_ASAP7_6t_L U453 ( .A(n42), .Y(n191) );
  XOR2xp5r_ASAP7_6t_L U454 ( .A(n192), .B(n193), .Y(n42) );
  XOR2xp5r_ASAP7_6t_L U455 ( .A(n188), .B(n187), .Y(n193) );
  OAI22xp5_ASAP7_6t_L U456 ( .A1(n194), .A2(n195), .B1(n196), .B2(n197), .Y(
        n187) );
  XOR2xp5r_ASAP7_6t_L U457 ( .A(n198), .B(n190), .Y(n197) );
  XOR2xp5r_ASAP7_6t_L U458 ( .A(n199), .B(n190), .Y(n195) );
  XOR2xp5r_ASAP7_6t_L U459 ( .A(n154), .B(n149), .Y(n190) );
  INVx1_ASAP7_6t_L U460 ( .A(n151), .Y(n149) );
  XOR2xp5r_ASAP7_6t_L U461 ( .A(n153), .B(n200), .Y(n151) );
  XOR2xp5r_ASAP7_6t_L U462 ( .A(n163), .B(n164), .Y(n200) );
  INVx1_ASAP7_6t_L U463 ( .A(n162), .Y(n164) );
  AOI22xp25_ASAP7_6t_L U464 ( .A1(n201), .A2(n202), .B1(n203), .B2(n204), .Y(
        n162) );
  XOR2xp5r_ASAP7_6t_L U465 ( .A(n205), .B(n165), .Y(n204) );
  XOR2xp5r_ASAP7_6t_L U466 ( .A(n206), .B(n165), .Y(n202) );
  XOR2xp5r_ASAP7_6t_L U467 ( .A(n207), .B(n208), .Y(n165) );
  XOR2xp5r_ASAP7_6t_L U468 ( .A(n160), .B(n158), .Y(n163) );
  AOI21xp25_ASAP7_6t_L U469 ( .A1(n209), .A2(n210), .B(n211), .Y(n158) );
  NOR3x1f_ASAP7_6t_L U470 ( .A(n210), .B(n212), .C(n213), .Y(n211) );
  INVx1_ASAP7_6t_L U471 ( .A(n159), .Y(n160) );
  XOR2xp5r_ASAP7_6t_L U472 ( .A(n214), .B(n215), .Y(n159) );
  XOR2xp5r_ASAP7_6t_L U473 ( .A(n216), .B(n161), .Y(n214) );
  NAND2xp5R_ASAP7_6t_L U474 ( .A(a[7]), .B(b[7]), .Y(n161) );
  NAND2xp5R_ASAP7_6t_L U475 ( .A(b[8]), .B(a[6]), .Y(n216) );
  AOI22xp25_ASAP7_6t_L U476 ( .A1(n217), .A2(n218), .B1(n219), .B2(n220), .Y(
        n153) );
  OA22x1_ASAP7_6t_L U477 ( .A1(n221), .A2(n222), .B1(n223), .B2(n224), .Y(n154) );
  INVx1_ASAP7_6t_L U478 ( .A(n196), .Y(n194) );
  XOR2xp5r_ASAP7_6t_L U479 ( .A(n185), .B(n184), .Y(n188) );
  XOR2xp5r_ASAP7_6t_L U480 ( .A(n167), .B(n225), .Y(n184) );
  XOR2xp5r_ASAP7_6t_L U481 ( .A(n226), .B(n166), .Y(n225) );
  XOR2xp5r_ASAP7_6t_L U482 ( .A(n227), .B(n169), .Y(n166) );
  XOR2xp5r_ASAP7_6t_L U483 ( .A(n171), .B(n176), .Y(n169) );
  AO21x1_ASAP7_6t_L U484 ( .A1(n228), .A2(n229), .B(n230), .Y(n176) );
  NOR3x1f_ASAP7_6t_L U485 ( .A(n229), .B(n231), .C(n232), .Y(n230) );
  XOR2xp5r_ASAP7_6t_L U486 ( .A(n233), .B(n234), .Y(n171) );
  XOR2xp5r_ASAP7_6t_L U487 ( .A(n175), .B(n235), .Y(n234) );
  NAND2xp5R_ASAP7_6t_L U488 ( .A(b[4]), .B(a[10]), .Y(n235) );
  NOR2xp5_ASAP7_6t_L U489 ( .A(n236), .B(n231), .Y(n175) );
  NOR2xp5_ASAP7_6t_L U490 ( .A(n237), .B(n238), .Y(n227) );
  NOR2xp5_ASAP7_6t_L U491 ( .A(n104), .B(n89), .Y(n226) );
  XOR2xp5r_ASAP7_6t_L U492 ( .A(n183), .B(n239), .Y(n167) );
  NAND2xp5R_ASAP7_6t_L U493 ( .A(b[1]), .B(a[13]), .Y(n239) );
  NAND2xp5R_ASAP7_6t_L U494 ( .A(b[2]), .B(a[12]), .Y(n183) );
  AO21x1_ASAP7_6t_L U495 ( .A1(n238), .A2(n240), .B(n241), .Y(n185) );
  NOR3x1f_ASAP7_6t_L U496 ( .A(n240), .B(n242), .C(n93), .Y(n241) );
  AOI22xp25_ASAP7_6t_L U497 ( .A1(n243), .A2(n244), .B1(n245), .B2(n246), .Y(
        n192) );
  OA22x1_ASAP7_6t_L U498 ( .A1(n247), .A2(n248), .B1(n249), .B2(n250), .Y(n41)
         );
  INVx1_ASAP7_6t_L U499 ( .A(n249), .Y(n247) );
  AO22x1_ASAP7_6t_L U500 ( .A1(n43), .A2(n44), .B1(n251), .B2(n252), .Y(c[95])
         );
  INVx1_ASAP7_6t_L U501 ( .A(n251), .Y(n44) );
  XOR2xp5r_ASAP7_6t_L U502 ( .A(n252), .B(n253), .Y(n251) );
  XOR2xp5r_ASAP7_6t_L U503 ( .A(n248), .B(n249), .Y(n253) );
  XOR2xp5r_ASAP7_6t_L U504 ( .A(n254), .B(n250), .Y(n249) );
  XOR2xp5r_ASAP7_6t_L U505 ( .A(n199), .B(n196), .Y(n250) );
  XOR2xp5r_ASAP7_6t_L U506 ( .A(n198), .B(n255), .Y(n196) );
  XOR2xp5r_ASAP7_6t_L U507 ( .A(n222), .B(n223), .Y(n255) );
  INVx1_ASAP7_6t_L U508 ( .A(n221), .Y(n223) );
  AOI22xp25_ASAP7_6t_L U509 ( .A1(n256), .A2(n257), .B1(n258), .B2(n259), .Y(
        n221) );
  XOR2xp5r_ASAP7_6t_L U510 ( .A(n260), .B(n224), .Y(n259) );
  XOR2xp5r_ASAP7_6t_L U511 ( .A(n261), .B(n224), .Y(n257) );
  XOR2xp5r_ASAP7_6t_L U512 ( .A(n201), .B(n206), .Y(n224) );
  AOI21xp25_ASAP7_6t_L U513 ( .A1(n262), .A2(n263), .B(n264), .Y(n206) );
  NOR3x1f_ASAP7_6t_L U514 ( .A(n263), .B(n265), .C(n90), .Y(n264) );
  INVx1_ASAP7_6t_L U515 ( .A(n203), .Y(n201) );
  XOR2xp5r_ASAP7_6t_L U516 ( .A(n266), .B(n267), .Y(n203) );
  XOR2xp5r_ASAP7_6t_L U517 ( .A(n205), .B(n268), .Y(n267) );
  NAND2xp5R_ASAP7_6t_L U518 ( .A(a[2]), .B(b[11]), .Y(n268) );
  NAND2xp5R_ASAP7_6t_L U519 ( .A(a[3]), .B(b[10]), .Y(n205) );
  XOR2xp5r_ASAP7_6t_L U520 ( .A(n219), .B(n217), .Y(n222) );
  AO21x1_ASAP7_6t_L U521 ( .A1(n269), .A2(n270), .B(n271), .Y(n217) );
  NOR3x1f_ASAP7_6t_L U522 ( .A(n270), .B(n272), .C(n213), .Y(n271) );
  INVx1_ASAP7_6t_L U523 ( .A(n218), .Y(n219) );
  XOR2xp5r_ASAP7_6t_L U524 ( .A(n210), .B(n273), .Y(n218) );
  XOR2xp5r_ASAP7_6t_L U525 ( .A(n220), .B(n274), .Y(n273) );
  NAND2xp5R_ASAP7_6t_L U526 ( .A(a[6]), .B(b[7]), .Y(n274) );
  NOR2xp5_ASAP7_6t_L U527 ( .A(n275), .B(n272), .Y(n220) );
  XOR2xp5r_ASAP7_6t_L U528 ( .A(n276), .B(n209), .Y(n210) );
  NOR2xp5_ASAP7_6t_L U529 ( .A(n277), .B(n278), .Y(n209) );
  NAND2xp5R_ASAP7_6t_L U530 ( .A(a[5]), .B(b[8]), .Y(n276) );
  AOI22xp25_ASAP7_6t_L U531 ( .A1(n279), .A2(n280), .B1(n281), .B2(n282), .Y(
        n198) );
  OA22x1_ASAP7_6t_L U532 ( .A1(n283), .A2(n284), .B1(n285), .B2(n286), .Y(n199) );
  INVx1_ASAP7_6t_L U533 ( .A(n283), .Y(n285) );
  AOI21xp25_ASAP7_6t_L U534 ( .A1(n287), .A2(n288), .B(n289), .Y(n254) );
  NOR3x1f_ASAP7_6t_L U535 ( .A(n287), .B(n290), .C(n291), .Y(n289) );
  INVx1_ASAP7_6t_L U536 ( .A(n292), .Y(n288) );
  XOR2xp5r_ASAP7_6t_L U537 ( .A(n243), .B(n245), .Y(n248) );
  INVx1_ASAP7_6t_L U538 ( .A(n244), .Y(n245) );
  XOR2xp5r_ASAP7_6t_L U539 ( .A(n240), .B(n293), .Y(n244) );
  XOR2xp5r_ASAP7_6t_L U540 ( .A(n246), .B(n294), .Y(n293) );
  NAND2xp5R_ASAP7_6t_L U541 ( .A(b[1]), .B(a[12]), .Y(n294) );
  NOR2xp5_ASAP7_6t_L U542 ( .A(n89), .B(n102), .Y(n246) );
  XOR2xp5r_ASAP7_6t_L U543 ( .A(n238), .B(n295), .Y(n240) );
  NAND2xp5R_ASAP7_6t_L U544 ( .A(n296), .B(n297), .Y(n295) );
  XOR2xp5r_ASAP7_6t_L U545 ( .A(n229), .B(n298), .Y(n238) );
  XOR2xp5r_ASAP7_6t_L U546 ( .A(n299), .B(n237), .Y(n298) );
  NAND2xp5R_ASAP7_6t_L U547 ( .A(a[11]), .B(b[2]), .Y(n237) );
  NOR2xp5_ASAP7_6t_L U548 ( .A(n231), .B(n232), .Y(n299) );
  XOR2xp5r_ASAP7_6t_L U549 ( .A(n300), .B(n228), .Y(n229) );
  NOR2xp5_ASAP7_6t_L U550 ( .A(n301), .B(n302), .Y(n228) );
  NAND2xp5R_ASAP7_6t_L U551 ( .A(a[9]), .B(b[4]), .Y(n300) );
  AO21x1_ASAP7_6t_L U552 ( .A1(n303), .A2(n304), .B(n305), .Y(n243) );
  NOR3x1f_ASAP7_6t_L U553 ( .A(n304), .B(n93), .C(n236), .Y(n305) );
  OAI22xp5_ASAP7_6t_L U554 ( .A1(n306), .A2(n307), .B1(n308), .B2(n309), .Y(
        n252) );
  OAI22xp5_ASAP7_6t_L U555 ( .A1(n310), .A2(n311), .B1(n312), .B2(n313), .Y(
        n43) );
  INVx1_ASAP7_6t_L U556 ( .A(n312), .Y(n310) );
  AO22x1_ASAP7_6t_L U557 ( .A1(n45), .A2(n46), .B1(n314), .B2(n315), .Y(c[94])
         );
  INVx1_ASAP7_6t_L U558 ( .A(n314), .Y(n46) );
  XOR2xp5r_ASAP7_6t_L U559 ( .A(n315), .B(n316), .Y(n314) );
  XOR2xp5r_ASAP7_6t_L U560 ( .A(n311), .B(n312), .Y(n316) );
  OAI22xp5_ASAP7_6t_L U561 ( .A1(n317), .A2(n318), .B1(n319), .B2(n320), .Y(
        n312) );
  XOR2xp5r_ASAP7_6t_L U562 ( .A(n321), .B(n313), .Y(n320) );
  INVx1_ASAP7_6t_L U563 ( .A(n322), .Y(n318) );
  XOR2xp5r_ASAP7_6t_L U564 ( .A(n323), .B(n313), .Y(n322) );
  XOR2xp5r_ASAP7_6t_L U565 ( .A(n292), .B(n287), .Y(n313) );
  XOR2xp5r_ASAP7_6t_L U566 ( .A(n324), .B(n283), .Y(n287) );
  AOI22xp25_ASAP7_6t_L U567 ( .A1(n325), .A2(n326), .B1(n327), .B2(n328), .Y(
        n283) );
  XOR2xp5r_ASAP7_6t_L U568 ( .A(n329), .B(n286), .Y(n328) );
  XOR2xp5r_ASAP7_6t_L U569 ( .A(n330), .B(n286), .Y(n326) );
  XOR2xp5r_ASAP7_6t_L U570 ( .A(n256), .B(n261), .Y(n286) );
  AOI21xp25_ASAP7_6t_L U571 ( .A1(n331), .A2(n332), .B(n333), .Y(n261) );
  NOR3x1f_ASAP7_6t_L U572 ( .A(n332), .B(n277), .C(n90), .Y(n333) );
  INVx1_ASAP7_6t_L U573 ( .A(n258), .Y(n256) );
  XOR2xp5r_ASAP7_6t_L U574 ( .A(n334), .B(n263), .Y(n258) );
  XOR2xp5r_ASAP7_6t_L U575 ( .A(n335), .B(n262), .Y(n263) );
  NOR2xp5_ASAP7_6t_L U576 ( .A(n336), .B(n94), .Y(n262) );
  NAND2xp5R_ASAP7_6t_L U577 ( .A(b[11]), .B(a[1]), .Y(n335) );
  XOR2xp5r_ASAP7_6t_L U578 ( .A(n337), .B(n260), .Y(n334) );
  NAND2xp5R_ASAP7_6t_L U579 ( .A(a[3]), .B(b[9]), .Y(n260) );
  NAND2xp5R_ASAP7_6t_L U580 ( .A(a[2]), .B(b[10]), .Y(n337) );
  INVx1_ASAP7_6t_L U581 ( .A(n327), .Y(n325) );
  XOR2xp5r_ASAP7_6t_L U582 ( .A(n338), .B(n284), .Y(n324) );
  XOR2xp5r_ASAP7_6t_L U583 ( .A(n281), .B(n279), .Y(n284) );
  AO21x1_ASAP7_6t_L U584 ( .A1(n339), .A2(n340), .B(n341), .Y(n279) );
  NOR3x1f_ASAP7_6t_L U585 ( .A(n340), .B(n302), .C(n213), .Y(n341) );
  INVx1_ASAP7_6t_L U586 ( .A(n342), .Y(n340) );
  INVx1_ASAP7_6t_L U587 ( .A(n280), .Y(n281) );
  XOR2xp5r_ASAP7_6t_L U588 ( .A(n343), .B(n270), .Y(n280) );
  XOR2xp5r_ASAP7_6t_L U589 ( .A(n344), .B(n269), .Y(n270) );
  NOR2xp5_ASAP7_6t_L U590 ( .A(n345), .B(n278), .Y(n269) );
  NAND2xp5R_ASAP7_6t_L U591 ( .A(b[7]), .B(a[5]), .Y(n344) );
  XOR2xp5r_ASAP7_6t_L U592 ( .A(n346), .B(n282), .Y(n343) );
  NOR2xp5_ASAP7_6t_L U593 ( .A(n275), .B(n302), .Y(n282) );
  NAND2xp5R_ASAP7_6t_L U594 ( .A(a[6]), .B(b[6]), .Y(n346) );
  NOR2xp5_ASAP7_6t_L U595 ( .A(n291), .B(n290), .Y(n338) );
  AOI22xp25_ASAP7_6t_L U596 ( .A1(n347), .A2(n290), .B1(n348), .B2(n349), .Y(
        n292) );
  INVx1_ASAP7_6t_L U597 ( .A(n348), .Y(n347) );
  XOR2xp5r_ASAP7_6t_L U598 ( .A(n308), .B(n306), .Y(n311) );
  AOI21xp25_ASAP7_6t_L U599 ( .A1(n350), .A2(n351), .B(n352), .Y(n306) );
  NOR3x1f_ASAP7_6t_L U600 ( .A(n351), .B(n93), .C(n232), .Y(n352) );
  INVx1_ASAP7_6t_L U601 ( .A(n307), .Y(n308) );
  XOR2xp5r_ASAP7_6t_L U602 ( .A(n353), .B(n304), .Y(n307) );
  XOR2xp5r_ASAP7_6t_L U603 ( .A(n303), .B(n354), .Y(n304) );
  NAND2xp5R_ASAP7_6t_L U604 ( .A(a[10]), .B(b[2]), .Y(n354) );
  XOR2xp5r_ASAP7_6t_L U605 ( .A(n297), .B(n296), .Y(n303) );
  NOR2xp5_ASAP7_6t_L U606 ( .A(n355), .B(n301), .Y(n296) );
  NOR2xp5_ASAP7_6t_L U607 ( .A(n356), .B(n231), .Y(n297) );
  XOR2xp5r_ASAP7_6t_L U608 ( .A(n357), .B(n309), .Y(n353) );
  NAND2xp5R_ASAP7_6t_L U609 ( .A(b[0]), .B(a[12]), .Y(n309) );
  NAND2xp5R_ASAP7_6t_L U610 ( .A(a[11]), .B(b[1]), .Y(n357) );
  OAI22xp5_ASAP7_6t_L U611 ( .A1(n358), .A2(n359), .B1(n360), .B2(n361), .Y(
        n315) );
  OAI22xp5_ASAP7_6t_L U612 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .Y(
        n45) );
  INVx1_ASAP7_6t_L U613 ( .A(n364), .Y(n362) );
  OAI22xp5_ASAP7_6t_L U614 ( .A1(n47), .A2(n48), .B1(n366), .B2(n367), .Y(
        c[93]) );
  INVx1_ASAP7_6t_L U615 ( .A(n366), .Y(n48) );
  XOR2xp5r_ASAP7_6t_L U616 ( .A(n367), .B(n368), .Y(n366) );
  XOR2xp5r_ASAP7_6t_L U617 ( .A(n363), .B(n364), .Y(n368) );
  XOR2xp5r_ASAP7_6t_L U618 ( .A(n369), .B(n365), .Y(n364) );
  XOR2xp5r_ASAP7_6t_L U619 ( .A(n319), .B(n323), .Y(n365) );
  AOI22xp25_ASAP7_6t_L U620 ( .A1(n370), .A2(n371), .B1(n372), .B2(n373), .Y(
        n323) );
  INVx1_ASAP7_6t_L U621 ( .A(n370), .Y(n372) );
  INVx1_ASAP7_6t_L U622 ( .A(n317), .Y(n319) );
  XOR2xp5r_ASAP7_6t_L U623 ( .A(n374), .B(n348), .Y(n317) );
  AOI22xp25_ASAP7_6t_L U624 ( .A1(n375), .A2(n376), .B1(n377), .B2(n378), .Y(
        n348) );
  XOR2xp5r_ASAP7_6t_L U625 ( .A(n379), .B(n349), .Y(n378) );
  INVx1_ASAP7_6t_L U626 ( .A(n375), .Y(n377) );
  XOR2xp5r_ASAP7_6t_L U627 ( .A(n380), .B(n349), .Y(n376) );
  XOR2xp5r_ASAP7_6t_L U628 ( .A(n327), .B(n330), .Y(n349) );
  AOI21xp25_ASAP7_6t_L U629 ( .A1(n381), .A2(n382), .B(n383), .Y(n330) );
  NOR3x1f_ASAP7_6t_L U630 ( .A(n382), .B(n345), .C(n90), .Y(n383) );
  XOR2xp5r_ASAP7_6t_L U631 ( .A(n384), .B(n332), .Y(n327) );
  XOR2xp5r_ASAP7_6t_L U632 ( .A(n385), .B(n331), .Y(n332) );
  NOR2xp5_ASAP7_6t_L U633 ( .A(n94), .B(n386), .Y(n331) );
  NAND2xp5R_ASAP7_6t_L U634 ( .A(b[10]), .B(a[1]), .Y(n385) );
  XOR2xp5r_ASAP7_6t_L U635 ( .A(n387), .B(n329), .Y(n384) );
  NAND2xp5R_ASAP7_6t_L U636 ( .A(a[3]), .B(b[8]), .Y(n329) );
  NAND2xp5R_ASAP7_6t_L U637 ( .A(a[2]), .B(b[9]), .Y(n387) );
  XOR2xp5r_ASAP7_6t_L U638 ( .A(n321), .B(n290), .Y(n374) );
  XOR2xp5r_ASAP7_6t_L U639 ( .A(n388), .B(n342), .Y(n290) );
  XOR2xp5r_ASAP7_6t_L U640 ( .A(n389), .B(n339), .Y(n342) );
  NOR2xp5_ASAP7_6t_L U641 ( .A(n278), .B(n212), .Y(n339) );
  NOR2xp5_ASAP7_6t_L U642 ( .A(n272), .B(n390), .Y(n389) );
  XOR2xp5r_ASAP7_6t_L U643 ( .A(n391), .B(n291), .Y(n388) );
  NAND2xp5R_ASAP7_6t_L U644 ( .A(a[7]), .B(b[4]), .Y(n291) );
  NAND2xp5R_ASAP7_6t_L U645 ( .A(a[6]), .B(b[5]), .Y(n391) );
  NOR3x1f_ASAP7_6t_L U646 ( .A(n392), .B(n302), .C(n390), .Y(n321) );
  AOI21xp25_ASAP7_6t_L U647 ( .A1(n393), .A2(n394), .B(n395), .Y(n369) );
  NOR3x1f_ASAP7_6t_L U648 ( .A(n393), .B(n355), .C(n213), .Y(n395) );
  XOR2xp5r_ASAP7_6t_L U649 ( .A(n360), .B(n358), .Y(n363) );
  AOI21xp25_ASAP7_6t_L U650 ( .A1(n396), .A2(n397), .B(n398), .Y(n358) );
  NOR3x1f_ASAP7_6t_L U651 ( .A(n397), .B(n93), .C(n356), .Y(n398) );
  INVx1_ASAP7_6t_L U652 ( .A(n359), .Y(n360) );
  XOR2xp5r_ASAP7_6t_L U653 ( .A(n399), .B(n351), .Y(n359) );
  XOR2xp5r_ASAP7_6t_L U654 ( .A(n400), .B(n350), .Y(n351) );
  NOR2xp5_ASAP7_6t_L U655 ( .A(n301), .B(n231), .Y(n350) );
  NAND2xp5R_ASAP7_6t_L U656 ( .A(b[2]), .B(a[9]), .Y(n400) );
  XOR2xp5r_ASAP7_6t_L U657 ( .A(n401), .B(n361), .Y(n399) );
  NAND2xp5R_ASAP7_6t_L U658 ( .A(a[11]), .B(b[0]), .Y(n361) );
  NAND2xp5R_ASAP7_6t_L U659 ( .A(a[10]), .B(b[1]), .Y(n401) );
  OA22x1_ASAP7_6t_L U660 ( .A1(n402), .A2(n403), .B1(n404), .B2(n405), .Y(n367) );
  INVx1_ASAP7_6t_L U661 ( .A(n403), .Y(n404) );
  AOI22xp25_ASAP7_6t_L U662 ( .A1(n406), .A2(n407), .B1(n408), .B2(n409), .Y(
        n47) );
  INVx1_ASAP7_6t_L U663 ( .A(n408), .Y(n406) );
  AO22x1_ASAP7_6t_L U664 ( .A1(n49), .A2(n50), .B1(n410), .B2(n411), .Y(c[92])
         );
  INVx1_ASAP7_6t_L U665 ( .A(n410), .Y(n50) );
  XOR2xp5r_ASAP7_6t_L U666 ( .A(n411), .B(n412), .Y(n410) );
  XOR2xp5r_ASAP7_6t_L U667 ( .A(n407), .B(n408), .Y(n412) );
  AOI22xp25_ASAP7_6t_L U668 ( .A1(n413), .A2(n414), .B1(n415), .B2(n416), .Y(
        n408) );
  XOR2xp5r_ASAP7_6t_L U669 ( .A(n417), .B(n409), .Y(n416) );
  XOR2xp5r_ASAP7_6t_L U670 ( .A(n418), .B(n409), .Y(n414) );
  XOR2xp5r_ASAP7_6t_L U671 ( .A(n394), .B(n393), .Y(n409) );
  XOR2xp5r_ASAP7_6t_L U672 ( .A(n371), .B(n419), .Y(n393) );
  XOR2xp5r_ASAP7_6t_L U673 ( .A(n420), .B(n370), .Y(n419) );
  XOR2xp5r_ASAP7_6t_L U674 ( .A(n421), .B(n373), .Y(n370) );
  XOR2xp5r_ASAP7_6t_L U675 ( .A(n375), .B(n380), .Y(n373) );
  AO21x1_ASAP7_6t_L U676 ( .A1(n422), .A2(n423), .B(n424), .Y(n380) );
  NOR3x1f_ASAP7_6t_L U677 ( .A(n423), .B(n212), .C(n90), .Y(n424) );
  XOR2xp5r_ASAP7_6t_L U678 ( .A(n425), .B(n382), .Y(n375) );
  XOR2xp5r_ASAP7_6t_L U679 ( .A(n426), .B(n381), .Y(n382) );
  NOR2xp5_ASAP7_6t_L U680 ( .A(n94), .B(n265), .Y(n381) );
  NAND2xp5R_ASAP7_6t_L U681 ( .A(b[9]), .B(a[1]), .Y(n426) );
  XOR2xp5r_ASAP7_6t_L U682 ( .A(n427), .B(n379), .Y(n425) );
  NOR2xp5_ASAP7_6t_L U683 ( .A(n428), .B(n212), .Y(n379) );
  NAND2xp5R_ASAP7_6t_L U684 ( .A(a[2]), .B(b[8]), .Y(n427) );
  NOR2xp5_ASAP7_6t_L U685 ( .A(n429), .B(n430), .Y(n421) );
  NOR2xp5_ASAP7_6t_L U686 ( .A(n355), .B(n213), .Y(n420) );
  XOR2xp5r_ASAP7_6t_L U687 ( .A(n392), .B(n431), .Y(n371) );
  NAND2xp5R_ASAP7_6t_L U688 ( .A(a[5]), .B(b[5]), .Y(n431) );
  NAND2xp5R_ASAP7_6t_L U689 ( .A(a[4]), .B(b[6]), .Y(n392) );
  AO21x1_ASAP7_6t_L U690 ( .A1(n430), .A2(n432), .B(n433), .Y(n394) );
  NOR3x1f_ASAP7_6t_L U691 ( .A(n432), .B(n302), .C(n278), .Y(n433) );
  INVx1_ASAP7_6t_L U692 ( .A(n415), .Y(n413) );
  XOR2xp5r_ASAP7_6t_L U693 ( .A(n403), .B(n402), .Y(n407) );
  AOI21xp25_ASAP7_6t_L U694 ( .A1(n434), .A2(n435), .B(n436), .Y(n402) );
  NOR3x1f_ASAP7_6t_L U695 ( .A(n435), .B(n93), .C(n301), .Y(n436) );
  XOR2xp5r_ASAP7_6t_L U696 ( .A(n437), .B(n397), .Y(n403) );
  XOR2xp5r_ASAP7_6t_L U697 ( .A(n438), .B(n396), .Y(n397) );
  NOR2xp5_ASAP7_6t_L U698 ( .A(n275), .B(n231), .Y(n396) );
  NAND2xp5R_ASAP7_6t_L U699 ( .A(b[2]), .B(a[8]), .Y(n438) );
  XOR2xp5r_ASAP7_6t_L U700 ( .A(n439), .B(n405), .Y(n437) );
  NAND2xp5R_ASAP7_6t_L U701 ( .A(a[10]), .B(b[0]), .Y(n405) );
  NAND2xp5R_ASAP7_6t_L U702 ( .A(a[9]), .B(b[1]), .Y(n439) );
  OAI22xp5_ASAP7_6t_L U703 ( .A1(n440), .A2(n441), .B1(n442), .B2(n443), .Y(
        n411) );
  OAI22xp5_ASAP7_6t_L U704 ( .A1(n444), .A2(n445), .B1(n446), .B2(n447), .Y(
        n49) );
  OAI22xp5_ASAP7_6t_L U705 ( .A1(n51), .A2(n52), .B1(n448), .B2(n449), .Y(
        c[91]) );
  INVx1_ASAP7_6t_L U706 ( .A(n448), .Y(n52) );
  XOR2xp5r_ASAP7_6t_L U707 ( .A(n449), .B(n450), .Y(n448) );
  XOR2xp5r_ASAP7_6t_L U708 ( .A(n445), .B(n446), .Y(n450) );
  INVx1_ASAP7_6t_L U709 ( .A(n444), .Y(n446) );
  AOI22xp25_ASAP7_6t_L U710 ( .A1(n451), .A2(n452), .B1(n453), .B2(n454), .Y(
        n444) );
  XOR2xp5r_ASAP7_6t_L U711 ( .A(n455), .B(n447), .Y(n454) );
  XOR2xp5r_ASAP7_6t_L U712 ( .A(n456), .B(n447), .Y(n452) );
  XOR2xp5r_ASAP7_6t_L U713 ( .A(n418), .B(n415), .Y(n447) );
  XOR2xp5r_ASAP7_6t_L U714 ( .A(n432), .B(n457), .Y(n415) );
  XOR2xp5r_ASAP7_6t_L U715 ( .A(n458), .B(n417), .Y(n457) );
  NOR2xp5_ASAP7_6t_L U716 ( .A(n390), .B(n355), .Y(n417) );
  NOR2xp5_ASAP7_6t_L U717 ( .A(n302), .B(n278), .Y(n458) );
  XOR2xp5r_ASAP7_6t_L U718 ( .A(n430), .B(n459), .Y(n432) );
  NAND2xp5R_ASAP7_6t_L U719 ( .A(n460), .B(n461), .Y(n459) );
  XOR2xp5r_ASAP7_6t_L U720 ( .A(n462), .B(n463), .Y(n430) );
  XOR2xp5r_ASAP7_6t_L U721 ( .A(n429), .B(n464), .Y(n463) );
  NAND2xp5R_ASAP7_6t_L U722 ( .A(a[2]), .B(b[7]), .Y(n464) );
  NAND2xp5R_ASAP7_6t_L U723 ( .A(a[3]), .B(b[6]), .Y(n429) );
  INVx1_ASAP7_6t_L U724 ( .A(n423), .Y(n462) );
  XOR2xp5r_ASAP7_6t_L U725 ( .A(n465), .B(n422), .Y(n423) );
  NOR2xp5_ASAP7_6t_L U726 ( .A(n94), .B(n277), .Y(n422) );
  NAND2xp5R_ASAP7_6t_L U727 ( .A(b[8]), .B(a[1]), .Y(n465) );
  AO21x1_ASAP7_6t_L U728 ( .A1(n466), .A2(n467), .B(n468), .Y(n418) );
  NOR3x1f_ASAP7_6t_L U729 ( .A(n467), .B(n302), .C(n428), .Y(n468) );
  XOR2xp5r_ASAP7_6t_L U730 ( .A(n442), .B(n440), .Y(n445) );
  AOI21xp25_ASAP7_6t_L U731 ( .A1(n469), .A2(n470), .B(n471), .Y(n440) );
  NOR3x1f_ASAP7_6t_L U732 ( .A(n470), .B(n93), .C(n275), .Y(n471) );
  INVx1_ASAP7_6t_L U733 ( .A(n441), .Y(n442) );
  XOR2xp5r_ASAP7_6t_L U734 ( .A(n472), .B(n435), .Y(n441) );
  XOR2xp5r_ASAP7_6t_L U735 ( .A(n473), .B(n434), .Y(n435) );
  NOR2xp5_ASAP7_6t_L U736 ( .A(n213), .B(n231), .Y(n434) );
  NAND2xp5R_ASAP7_6t_L U737 ( .A(b[2]), .B(a[7]), .Y(n473) );
  XOR2xp5r_ASAP7_6t_L U738 ( .A(n474), .B(n443), .Y(n472) );
  NAND2xp5R_ASAP7_6t_L U739 ( .A(a[9]), .B(b[0]), .Y(n443) );
  NAND2xp5R_ASAP7_6t_L U740 ( .A(a[8]), .B(b[1]), .Y(n474) );
  AOI22xp25_ASAP7_6t_L U741 ( .A1(n475), .A2(n476), .B1(n477), .B2(n478), .Y(
        n449) );
  OA22x1_ASAP7_6t_L U742 ( .A1(n479), .A2(n480), .B1(n481), .B2(n482), .Y(n51)
         );
  INVx1_ASAP7_6t_L U743 ( .A(n479), .Y(n481) );
  AO21x1_ASAP7_6t_L U744 ( .A1(n54), .A2(n53), .B(n483), .Y(c[90]) );
  NOR3x1f_ASAP7_6t_L U745 ( .A(n54), .B(n484), .C(n485), .Y(n483) );
  OAI22xp5_ASAP7_6t_L U746 ( .A1(n486), .A2(n487), .B1(n488), .B2(n489), .Y(
        n53) );
  XOR2xp5r_ASAP7_6t_L U747 ( .A(n490), .B(n479), .Y(n54) );
  AOI22xp25_ASAP7_6t_L U748 ( .A1(n491), .A2(n492), .B1(n493), .B2(n494), .Y(
        n479) );
  XOR2xp5r_ASAP7_6t_L U749 ( .A(n495), .B(n482), .Y(n494) );
  XOR2xp5r_ASAP7_6t_L U750 ( .A(n496), .B(n482), .Y(n492) );
  XOR2xp5r_ASAP7_6t_L U751 ( .A(n451), .B(n456), .Y(n482) );
  AOI21xp25_ASAP7_6t_L U752 ( .A1(n497), .A2(n498), .B(n499), .Y(n456) );
  NOR3x1f_ASAP7_6t_L U753 ( .A(n498), .B(n302), .C(n90), .Y(n499) );
  INVx1_ASAP7_6t_L U754 ( .A(n453), .Y(n451) );
  XOR2xp5r_ASAP7_6t_L U755 ( .A(n500), .B(n467), .Y(n453) );
  XOR2xp5r_ASAP7_6t_L U756 ( .A(n466), .B(n501), .Y(n467) );
  NAND2xp5R_ASAP7_6t_L U757 ( .A(a[2]), .B(b[6]), .Y(n501) );
  XOR2xp5r_ASAP7_6t_L U758 ( .A(n461), .B(n460), .Y(n466) );
  NOR2xp5_ASAP7_6t_L U759 ( .A(n94), .B(n345), .Y(n460) );
  NOR2xp5_ASAP7_6t_L U760 ( .A(n95), .B(n212), .Y(n461) );
  XOR2xp5r_ASAP7_6t_L U761 ( .A(n502), .B(n455), .Y(n500) );
  NAND2xp5R_ASAP7_6t_L U762 ( .A(a[4]), .B(b[4]), .Y(n455) );
  NAND2xp5R_ASAP7_6t_L U763 ( .A(a[3]), .B(b[5]), .Y(n502) );
  XOR2xp5r_ASAP7_6t_L U764 ( .A(n503), .B(n480), .Y(n490) );
  XOR2xp5r_ASAP7_6t_L U765 ( .A(n477), .B(n475), .Y(n480) );
  AO21x1_ASAP7_6t_L U766 ( .A1(n504), .A2(n505), .B(n506), .Y(n475) );
  NOR3x1f_ASAP7_6t_L U767 ( .A(n505), .B(n93), .C(n213), .Y(n506) );
  INVx1_ASAP7_6t_L U768 ( .A(n476), .Y(n477) );
  XOR2xp5r_ASAP7_6t_L U769 ( .A(n470), .B(n507), .Y(n476) );
  XOR2xp5r_ASAP7_6t_L U770 ( .A(n478), .B(n508), .Y(n507) );
  NAND2xp5R_ASAP7_6t_L U771 ( .A(a[7]), .B(b[1]), .Y(n508) );
  NOR2xp5_ASAP7_6t_L U772 ( .A(n301), .B(n89), .Y(n478) );
  XOR2xp5r_ASAP7_6t_L U773 ( .A(n469), .B(n509), .Y(n470) );
  NAND2xp5R_ASAP7_6t_L U774 ( .A(a[6]), .B(b[2]), .Y(n509) );
  NOR2xp5_ASAP7_6t_L U775 ( .A(n390), .B(n231), .Y(n469) );
  NOR2xp5_ASAP7_6t_L U776 ( .A(n485), .B(n484), .Y(n503) );
  OAI22xp5_ASAP7_6t_L U777 ( .A1(n56), .A2(n55), .B1(n510), .B2(n511), .Y(
        c[89]) );
  INVx1_ASAP7_6t_L U778 ( .A(n512), .Y(n511) );
  INVx1_ASAP7_6t_L U779 ( .A(n55), .Y(n510) );
  XOR2xp5r_ASAP7_6t_L U780 ( .A(n513), .B(n486), .Y(n55) );
  INVx1_ASAP7_6t_L U781 ( .A(n488), .Y(n486) );
  OAI22xp5_ASAP7_6t_L U782 ( .A1(n514), .A2(n515), .B1(n516), .B2(n517), .Y(
        n488) );
  XOR2xp5r_ASAP7_6t_L U783 ( .A(n518), .B(n489), .Y(n517) );
  XOR2xp5r_ASAP7_6t_L U784 ( .A(n519), .B(n489), .Y(n515) );
  XOR2xp5r_ASAP7_6t_L U785 ( .A(n491), .B(n496), .Y(n489) );
  AOI21xp25_ASAP7_6t_L U786 ( .A1(n520), .A2(n521), .B(n522), .Y(n496) );
  NOR3x1f_ASAP7_6t_L U787 ( .A(n521), .B(n355), .C(n90), .Y(n522) );
  INVx1_ASAP7_6t_L U788 ( .A(n493), .Y(n491) );
  XOR2xp5r_ASAP7_6t_L U789 ( .A(n523), .B(n498), .Y(n493) );
  XOR2xp5r_ASAP7_6t_L U790 ( .A(n524), .B(n497), .Y(n498) );
  NOR2xp5_ASAP7_6t_L U791 ( .A(n94), .B(n212), .Y(n497) );
  NAND2xp5R_ASAP7_6t_L U792 ( .A(b[6]), .B(a[1]), .Y(n524) );
  XOR2xp5r_ASAP7_6t_L U793 ( .A(n525), .B(n495), .Y(n523) );
  NAND2xp5R_ASAP7_6t_L U794 ( .A(a[3]), .B(b[4]), .Y(n495) );
  NAND2xp5R_ASAP7_6t_L U795 ( .A(a[2]), .B(b[5]), .Y(n525) );
  INVx1_ASAP7_6t_L U796 ( .A(n516), .Y(n514) );
  XOR2xp5r_ASAP7_6t_L U797 ( .A(n512), .B(n484), .Y(n513) );
  INVx1_ASAP7_6t_L U798 ( .A(n487), .Y(n484) );
  XOR2xp5r_ASAP7_6t_L U799 ( .A(n505), .B(n526), .Y(n487) );
  XOR2xp5r_ASAP7_6t_L U800 ( .A(n485), .B(n527), .Y(n526) );
  NAND2xp5R_ASAP7_6t_L U801 ( .A(a[6]), .B(b[1]), .Y(n527) );
  NAND2xp5R_ASAP7_6t_L U802 ( .A(a[7]), .B(b[0]), .Y(n485) );
  XOR2xp5r_ASAP7_6t_L U803 ( .A(n528), .B(n504), .Y(n505) );
  NOR2xp5_ASAP7_6t_L U804 ( .A(n278), .B(n231), .Y(n504) );
  NAND2xp5R_ASAP7_6t_L U805 ( .A(b[2]), .B(a[5]), .Y(n528) );
  NOR3x1f_ASAP7_6t_L U806 ( .A(n529), .B(n93), .C(n390), .Y(n512) );
  AOI22xp25_ASAP7_6t_L U807 ( .A1(n530), .A2(n531), .B1(n532), .B2(n533), .Y(
        n56) );
  INVx1_ASAP7_6t_L U808 ( .A(n530), .Y(n532) );
  AO21x1_ASAP7_6t_L U809 ( .A1(n58), .A2(n57), .B(n534), .Y(c[88]) );
  NOR3x1f_ASAP7_6t_L U810 ( .A(n58), .B(n89), .C(n213), .Y(n534) );
  AO21x1_ASAP7_6t_L U811 ( .A1(n535), .A2(n536), .B(n537), .Y(n57) );
  NOR3x1f_ASAP7_6t_L U812 ( .A(n536), .B(n93), .C(n278), .Y(n537) );
  XOR2xp5r_ASAP7_6t_L U813 ( .A(n531), .B(n538), .Y(n58) );
  XOR2xp5r_ASAP7_6t_L U814 ( .A(n539), .B(n530), .Y(n538) );
  XOR2xp5r_ASAP7_6t_L U815 ( .A(n540), .B(n533), .Y(n530) );
  XOR2xp5r_ASAP7_6t_L U816 ( .A(n516), .B(n519), .Y(n533) );
  AO21x1_ASAP7_6t_L U817 ( .A1(n541), .A2(n542), .B(n543), .Y(n519) );
  NOR3x1f_ASAP7_6t_L U818 ( .A(n542), .B(n231), .C(n90), .Y(n543) );
  XOR2xp5r_ASAP7_6t_L U819 ( .A(n521), .B(n544), .Y(n516) );
  XOR2xp5r_ASAP7_6t_L U820 ( .A(n518), .B(n545), .Y(n544) );
  NAND2xp5R_ASAP7_6t_L U821 ( .A(a[2]), .B(b[4]), .Y(n545) );
  NOR2xp5_ASAP7_6t_L U822 ( .A(n428), .B(n231), .Y(n518) );
  XOR2xp5r_ASAP7_6t_L U823 ( .A(n520), .B(n546), .Y(n521) );
  NAND2xp5R_ASAP7_6t_L U824 ( .A(a[1]), .B(b[5]), .Y(n546) );
  NOR2xp5_ASAP7_6t_L U825 ( .A(n94), .B(n272), .Y(n520) );
  NOR2xp5_ASAP7_6t_L U826 ( .A(n547), .B(n535), .Y(n540) );
  NOR2xp5_ASAP7_6t_L U827 ( .A(n89), .B(n213), .Y(n539) );
  INVx1_ASAP7_6t_L U828 ( .A(b[0]), .Y(n89) );
  XOR2xp5r_ASAP7_6t_L U829 ( .A(n529), .B(n548), .Y(n531) );
  NAND2xp5R_ASAP7_6t_L U830 ( .A(a[5]), .B(b[1]), .Y(n548) );
  NAND2xp5R_ASAP7_6t_L U831 ( .A(a[4]), .B(b[2]), .Y(n529) );
  OAI22xp5_ASAP7_6t_L U832 ( .A1(n59), .A2(n60), .B1(n549), .B2(n550), .Y(
        c[87]) );
  INVx1_ASAP7_6t_L U833 ( .A(n60), .Y(n549) );
  XOR2xp5r_ASAP7_6t_L U834 ( .A(n536), .B(n551), .Y(n60) );
  XOR2xp5r_ASAP7_6t_L U835 ( .A(n550), .B(n552), .Y(n551) );
  NAND2xp5R_ASAP7_6t_L U836 ( .A(a[4]), .B(b[1]), .Y(n552) );
  NAND2xp5R_ASAP7_6t_L U837 ( .A(a[5]), .B(b[0]), .Y(n550) );
  XOR2xp5r_ASAP7_6t_L U838 ( .A(n535), .B(n553), .Y(n536) );
  NAND2xp5R_ASAP7_6t_L U839 ( .A(n554), .B(n555), .Y(n553) );
  XOR2xp5r_ASAP7_6t_L U840 ( .A(n556), .B(n557), .Y(n535) );
  XOR2xp5r_ASAP7_6t_L U841 ( .A(n547), .B(n558), .Y(n557) );
  NAND2xp5R_ASAP7_6t_L U842 ( .A(a[2]), .B(b[3]), .Y(n558) );
  NAND2xp5R_ASAP7_6t_L U843 ( .A(a[3]), .B(b[2]), .Y(n547) );
  INVx1_ASAP7_6t_L U844 ( .A(n542), .Y(n556) );
  XOR2xp5r_ASAP7_6t_L U845 ( .A(n559), .B(n541), .Y(n542) );
  NOR2xp5_ASAP7_6t_L U846 ( .A(n94), .B(n302), .Y(n541) );
  NAND2xp5R_ASAP7_6t_L U847 ( .A(b[4]), .B(a[1]), .Y(n559) );
  AOI21xp25_ASAP7_6t_L U848 ( .A1(n560), .A2(n561), .B(n562), .Y(n59) );
  NOR3x1f_ASAP7_6t_L U849 ( .A(n561), .B(n93), .C(n428), .Y(n562) );
  OAI22xp5_ASAP7_6t_L U850 ( .A1(n62), .A2(n61), .B1(n563), .B2(n564), .Y(
        c[86]) );
  INVx1_ASAP7_6t_L U851 ( .A(n61), .Y(n563) );
  XOR2xp5r_ASAP7_6t_L U852 ( .A(n565), .B(n561), .Y(n61) );
  XOR2xp5r_ASAP7_6t_L U853 ( .A(n560), .B(n566), .Y(n561) );
  NAND2xp5R_ASAP7_6t_L U854 ( .A(a[2]), .B(b[2]), .Y(n566) );
  XOR2xp5r_ASAP7_6t_L U855 ( .A(n555), .B(n554), .Y(n560) );
  NOR2xp5_ASAP7_6t_L U856 ( .A(n94), .B(n355), .Y(n554) );
  NOR2xp5_ASAP7_6t_L U857 ( .A(n95), .B(n231), .Y(n555) );
  XOR2xp5r_ASAP7_6t_L U858 ( .A(n567), .B(n564), .Y(n565) );
  NAND2xp5R_ASAP7_6t_L U859 ( .A(a[4]), .B(b[0]), .Y(n564) );
  NAND2xp5R_ASAP7_6t_L U860 ( .A(a[3]), .B(b[1]), .Y(n567) );
  AOI21xp25_ASAP7_6t_L U861 ( .A1(n568), .A2(n569), .B(n570), .Y(n62) );
  NOR3x1f_ASAP7_6t_L U862 ( .A(n569), .B(n93), .C(n90), .Y(n570) );
  INVx1_ASAP7_6t_L U863 ( .A(n571), .Y(n569) );
  NOR2xp5_ASAP7_6t_L U864 ( .A(n1173), .B(n572), .Y(c[85]) );
  XOR2xp5r_ASAP7_6t_L U865 ( .A(n573), .B(n571), .Y(n1173) );
  XOR2xp5r_ASAP7_6t_L U866 ( .A(n574), .B(n568), .Y(n571) );
  NOR2xp5_ASAP7_6t_L U867 ( .A(n94), .B(n231), .Y(n568) );
  AND2x2_ASAP7_6t_L U868 ( .A(b[2]), .B(a[1]), .Y(n574) );
  XOR2xp5r_ASAP7_6t_L U869 ( .A(n575), .B(n572), .Y(n573) );
  NAND2xp5R_ASAP7_6t_L U870 ( .A(a[3]), .B(b[0]), .Y(n572) );
  NAND2xp5R_ASAP7_6t_L U871 ( .A(a[2]), .B(b[1]), .Y(n575) );
  NOR3x1f_ASAP7_6t_L U872 ( .A(n64), .B(n93), .C(n95), .Y(c[84]) );
  NAND2xp5R_ASAP7_6t_L U873 ( .A(a[0]), .B(b[2]), .Y(n64) );
  OAI22xp5_ASAP7_6t_L U874 ( .A1(n576), .A2(n577), .B1(n67), .B2(n68), .Y(
        c[110]) );
  AOI21xp25_ASAP7_6t_L U875 ( .A1(n578), .A2(n579), .B(n580), .Y(n68) );
  NOR3x1f_ASAP7_6t_L U876 ( .A(n579), .B(n104), .C(n581), .Y(n580) );
  INVx1_ASAP7_6t_L U877 ( .A(n67), .Y(n576) );
  XOR2xp5r_ASAP7_6t_L U878 ( .A(n582), .B(n103), .Y(n67) );
  INVx1_ASAP7_6t_L U879 ( .A(n101), .Y(n103) );
  XOR2xp5r_ASAP7_6t_L U880 ( .A(n583), .B(n584), .Y(n101) );
  NAND2xp5R_ASAP7_6t_L U881 ( .A(b[15]), .B(a[13]), .Y(n584) );
  AOI22xp25_ASAP7_6t_L U882 ( .A1(n585), .A2(n586), .B1(n587), .B2(n588), .Y(
        n583) );
  XOR2xp5r_ASAP7_6t_L U883 ( .A(n589), .B(n577), .Y(n582) );
  NAND2xp5R_ASAP7_6t_L U884 ( .A(b[13]), .B(a[15]), .Y(n577) );
  NAND2xp5R_ASAP7_6t_L U885 ( .A(b[14]), .B(a[14]), .Y(n589) );
  OAI22xp5_ASAP7_6t_L U886 ( .A1(n70), .A2(n69), .B1(n590), .B2(n591), .Y(
        c[109]) );
  INVx1_ASAP7_6t_L U887 ( .A(n69), .Y(n590) );
  XOR2xp5r_ASAP7_6t_L U888 ( .A(n592), .B(n579), .Y(n69) );
  AOI22xp25_ASAP7_6t_L U889 ( .A1(n593), .A2(n594), .B1(n595), .B2(n596), .Y(
        n579) );
  XOR2xp5r_ASAP7_6t_L U890 ( .A(n597), .B(n578), .Y(n596) );
  INVx1_ASAP7_6t_L U891 ( .A(n593), .Y(n595) );
  XOR2xp5r_ASAP7_6t_L U892 ( .A(n598), .B(n578), .Y(n594) );
  XOR2xp5r_ASAP7_6t_L U893 ( .A(n588), .B(n587), .Y(n578) );
  AO21x1_ASAP7_6t_L U894 ( .A1(n599), .A2(n600), .B(n601), .Y(n587) );
  NOR3x1f_ASAP7_6t_L U895 ( .A(n600), .B(n102), .C(n581), .Y(n601) );
  XOR2xp5r_ASAP7_6t_L U896 ( .A(n586), .B(n585), .Y(n588) );
  NOR2xp5_ASAP7_6t_L U897 ( .A(n98), .B(n102), .Y(n585) );
  NOR2xp5_ASAP7_6t_L U898 ( .A(n92), .B(n242), .Y(n586) );
  XOR2xp5r_ASAP7_6t_L U899 ( .A(n602), .B(n591), .Y(n592) );
  NAND2xp5R_ASAP7_6t_L U900 ( .A(b[12]), .B(a[15]), .Y(n591) );
  NAND2xp5R_ASAP7_6t_L U901 ( .A(b[13]), .B(a[14]), .Y(n602) );
  AOI21xp25_ASAP7_6t_L U902 ( .A1(n603), .A2(n604), .B(n605), .Y(n70) );
  NOR3x1f_ASAP7_6t_L U903 ( .A(n604), .B(n91), .C(n386), .Y(n605) );
  AO22x1_ASAP7_6t_L U904 ( .A1(n606), .A2(n607), .B1(n72), .B2(n71), .Y(c[108]) );
  OAI22xp5_ASAP7_6t_L U905 ( .A1(n608), .A2(n609), .B1(n610), .B2(n611), .Y(
        n71) );
  INVx1_ASAP7_6t_L U906 ( .A(n610), .Y(n608) );
  INVx1_ASAP7_6t_L U907 ( .A(n72), .Y(n607) );
  XOR2xp5r_ASAP7_6t_L U908 ( .A(n612), .B(n604), .Y(n72) );
  AOI22xp25_ASAP7_6t_L U909 ( .A1(n613), .A2(n614), .B1(n615), .B2(n616), .Y(
        n604) );
  XOR2xp5r_ASAP7_6t_L U910 ( .A(n617), .B(n603), .Y(n616) );
  XOR2xp5r_ASAP7_6t_L U911 ( .A(n618), .B(n603), .Y(n614) );
  XOR2xp5r_ASAP7_6t_L U912 ( .A(n593), .B(n598), .Y(n603) );
  AO21x1_ASAP7_6t_L U913 ( .A1(n619), .A2(n620), .B(n621), .Y(n598) );
  NOR3x1f_ASAP7_6t_L U914 ( .A(n620), .B(n242), .C(n581), .Y(n621) );
  XOR2xp5r_ASAP7_6t_L U915 ( .A(n622), .B(n600), .Y(n593) );
  XOR2xp5r_ASAP7_6t_L U916 ( .A(n623), .B(n599), .Y(n600) );
  NOR2xp5_ASAP7_6t_L U917 ( .A(n92), .B(n236), .Y(n599) );
  NAND2xp5R_ASAP7_6t_L U918 ( .A(a[12]), .B(b[14]), .Y(n623) );
  XOR2xp5r_ASAP7_6t_L U919 ( .A(n624), .B(n597), .Y(n622) );
  NOR2xp5_ASAP7_6t_L U920 ( .A(n336), .B(n104), .Y(n597) );
  NAND2xp5R_ASAP7_6t_L U921 ( .A(b[13]), .B(a[13]), .Y(n624) );
  XOR2xp5r_ASAP7_6t_L U922 ( .A(n625), .B(n606), .Y(n612) );
  NAND2xp5R_ASAP7_6t_L U923 ( .A(b[11]), .B(a[15]), .Y(n625) );
  OAI22xp5_ASAP7_6t_L U924 ( .A1(n626), .A2(n627), .B1(n628), .B2(n629), .Y(
        n606) );
  INVx1_ASAP7_6t_L U925 ( .A(n630), .Y(n627) );
  OAI22xp5_ASAP7_6t_L U926 ( .A1(n74), .A2(n73), .B1(n631), .B2(n632), .Y(
        c[107]) );
  INVx1_ASAP7_6t_L U927 ( .A(n631), .Y(n73) );
  XOR2xp5r_ASAP7_6t_L U928 ( .A(n632), .B(n633), .Y(n631) );
  XOR2xp5r_ASAP7_6t_L U929 ( .A(n609), .B(n610), .Y(n633) );
  OAI22xp5_ASAP7_6t_L U930 ( .A1(n634), .A2(n635), .B1(n636), .B2(n637), .Y(
        n610) );
  XOR2xp5r_ASAP7_6t_L U931 ( .A(n611), .B(n638), .Y(n637) );
  XOR2xp5r_ASAP7_6t_L U932 ( .A(n639), .B(n611), .Y(n635) );
  XOR2xp5r_ASAP7_6t_L U933 ( .A(n618), .B(n615), .Y(n611) );
  INVx1_ASAP7_6t_L U934 ( .A(n613), .Y(n615) );
  XOR2xp5r_ASAP7_6t_L U935 ( .A(n640), .B(n620), .Y(n613) );
  XOR2xp5r_ASAP7_6t_L U936 ( .A(n641), .B(n619), .Y(n620) );
  NOR2xp5_ASAP7_6t_L U937 ( .A(n92), .B(n232), .Y(n619) );
  NAND2xp5R_ASAP7_6t_L U938 ( .A(a[11]), .B(b[14]), .Y(n641) );
  XOR2xp5r_ASAP7_6t_L U939 ( .A(n642), .B(n617), .Y(n640) );
  NOR2xp5_ASAP7_6t_L U940 ( .A(n336), .B(n102), .Y(n617) );
  NAND2xp5R_ASAP7_6t_L U941 ( .A(b[13]), .B(a[12]), .Y(n642) );
  OR2x2_ASAP7_6t_L U942 ( .A(n643), .B(n644), .Y(n618) );
  NOR3x1f_ASAP7_6t_L U943 ( .A(n645), .B(n356), .C(n92), .Y(n644) );
  NOR3x1f_ASAP7_6t_L U944 ( .A(n646), .B(n232), .C(n98), .Y(n643) );
  INVx1_ASAP7_6t_L U945 ( .A(n645), .Y(n646) );
  INVx1_ASAP7_6t_L U946 ( .A(n636), .Y(n634) );
  XOR2xp5r_ASAP7_6t_L U947 ( .A(n630), .B(n626), .Y(n609) );
  AOI21xp25_ASAP7_6t_L U948 ( .A1(n647), .A2(n648), .B(n649), .Y(n626) );
  NOR3x1f_ASAP7_6t_L U949 ( .A(n648), .B(n104), .C(n265), .Y(n649) );
  XOR2xp5r_ASAP7_6t_L U950 ( .A(n628), .B(n629), .Y(n630) );
  NAND2xp5R_ASAP7_6t_L U951 ( .A(b[11]), .B(a[14]), .Y(n629) );
  NAND2xp5R_ASAP7_6t_L U952 ( .A(b[10]), .B(a[15]), .Y(n628) );
  AOI22xp25_ASAP7_6t_L U953 ( .A1(n650), .A2(n651), .B1(n652), .B2(n653), .Y(
        n632) );
  OA22x1_ASAP7_6t_L U954 ( .A1(n654), .A2(n655), .B1(n656), .B2(n657), .Y(n74)
         );
  OAI22xp5_ASAP7_6t_L U955 ( .A1(n76), .A2(n75), .B1(n658), .B2(n659), .Y(
        c[106]) );
  INVx1_ASAP7_6t_L U956 ( .A(n658), .Y(n75) );
  XOR2xp5r_ASAP7_6t_L U957 ( .A(n659), .B(n660), .Y(n658) );
  XOR2xp5r_ASAP7_6t_L U958 ( .A(n657), .B(n655), .Y(n660) );
  INVx1_ASAP7_6t_L U959 ( .A(n656), .Y(n655) );
  AOI22xp25_ASAP7_6t_L U960 ( .A1(n661), .A2(n662), .B1(n663), .B2(n664), .Y(
        n656) );
  XOR2xp5r_ASAP7_6t_L U961 ( .A(n665), .B(n654), .Y(n663) );
  XOR2xp5r_ASAP7_6t_L U962 ( .A(n666), .B(n654), .Y(n662) );
  XOR2xp5r_ASAP7_6t_L U963 ( .A(n636), .B(n638), .Y(n654) );
  AO21x1_ASAP7_6t_L U964 ( .A1(n667), .A2(n668), .B(n669), .Y(n638) );
  NOR3x1f_ASAP7_6t_L U965 ( .A(n668), .B(n232), .C(n581), .Y(n669) );
  XOR2xp5r_ASAP7_6t_L U966 ( .A(n670), .B(n645), .Y(n636) );
  XOR2xp5r_ASAP7_6t_L U967 ( .A(n671), .B(n672), .Y(n645) );
  NAND2xp5R_ASAP7_6t_L U968 ( .A(b[15]), .B(a[9]), .Y(n672) );
  AOI22xp25_ASAP7_6t_L U969 ( .A1(n673), .A2(n674), .B1(n675), .B2(n676), .Y(
        n671) );
  XOR2xp5r_ASAP7_6t_L U970 ( .A(n677), .B(n639), .Y(n670) );
  NOR2xp5_ASAP7_6t_L U971 ( .A(n581), .B(n236), .Y(n639) );
  NAND2xp5R_ASAP7_6t_L U972 ( .A(b[14]), .B(a[10]), .Y(n677) );
  XOR2xp5r_ASAP7_6t_L U973 ( .A(n652), .B(n650), .Y(n657) );
  AO21x1_ASAP7_6t_L U974 ( .A1(n678), .A2(n679), .B(n680), .Y(n650) );
  NOR3x1f_ASAP7_6t_L U975 ( .A(n679), .B(n104), .C(n277), .Y(n680) );
  INVx1_ASAP7_6t_L U976 ( .A(n651), .Y(n652) );
  XOR2xp5r_ASAP7_6t_L U977 ( .A(n648), .B(n681), .Y(n651) );
  XOR2xp5r_ASAP7_6t_L U978 ( .A(n653), .B(n682), .Y(n681) );
  NAND2xp5R_ASAP7_6t_L U979 ( .A(b[10]), .B(a[14]), .Y(n682) );
  NOR2xp5_ASAP7_6t_L U980 ( .A(n277), .B(n91), .Y(n653) );
  XOR2xp5r_ASAP7_6t_L U981 ( .A(n683), .B(n647), .Y(n648) );
  NOR2xp5_ASAP7_6t_L U982 ( .A(n336), .B(n242), .Y(n647) );
  NAND2xp5R_ASAP7_6t_L U983 ( .A(a[13]), .B(b[11]), .Y(n683) );
  AOI22xp25_ASAP7_6t_L U984 ( .A1(n684), .A2(n685), .B1(n686), .B2(n687), .Y(
        n659) );
  OA22x1_ASAP7_6t_L U985 ( .A1(n688), .A2(n689), .B1(n690), .B2(n691), .Y(n76)
         );
  OAI22xp5_ASAP7_6t_L U986 ( .A1(n78), .A2(n77), .B1(n692), .B2(n693), .Y(
        c[105]) );
  INVx1_ASAP7_6t_L U987 ( .A(n692), .Y(n77) );
  XOR2xp5r_ASAP7_6t_L U988 ( .A(n693), .B(n694), .Y(n692) );
  XOR2xp5r_ASAP7_6t_L U989 ( .A(n689), .B(n690), .Y(n694) );
  INVx1_ASAP7_6t_L U990 ( .A(n688), .Y(n690) );
  AOI22xp25_ASAP7_6t_L U991 ( .A1(n695), .A2(n696), .B1(n697), .B2(n698), .Y(
        n688) );
  XOR2xp5r_ASAP7_6t_L U992 ( .A(n699), .B(n691), .Y(n697) );
  XOR2xp5r_ASAP7_6t_L U993 ( .A(n700), .B(n691), .Y(n696) );
  XOR2xp5r_ASAP7_6t_L U994 ( .A(n664), .B(n665), .Y(n691) );
  AOI21xp25_ASAP7_6t_L U995 ( .A1(n701), .A2(n702), .B(n703), .Y(n665) );
  NOR3x1f_ASAP7_6t_L U996 ( .A(n702), .B(n236), .C(n386), .Y(n703) );
  INVx1_ASAP7_6t_L U997 ( .A(n661), .Y(n664) );
  XOR2xp5r_ASAP7_6t_L U998 ( .A(n704), .B(n668), .Y(n661) );
  AOI22xp25_ASAP7_6t_L U999 ( .A1(n705), .A2(n706), .B1(n707), .B2(n708), .Y(
        n668) );
  XOR2xp5r_ASAP7_6t_L U1000 ( .A(n709), .B(n667), .Y(n708) );
  INVx1_ASAP7_6t_L U1001 ( .A(n705), .Y(n707) );
  XOR2xp5r_ASAP7_6t_L U1002 ( .A(n710), .B(n667), .Y(n706) );
  XOR2xp5r_ASAP7_6t_L U1003 ( .A(n676), .B(n675), .Y(n667) );
  AO21x1_ASAP7_6t_L U1004 ( .A1(n711), .A2(n712), .B(n713), .Y(n675) );
  NOR3x1f_ASAP7_6t_L U1005 ( .A(n712), .B(n356), .C(n581), .Y(n713) );
  XOR2xp5r_ASAP7_6t_L U1006 ( .A(n674), .B(n673), .Y(n676) );
  NOR2xp5_ASAP7_6t_L U1007 ( .A(n98), .B(n356), .Y(n673) );
  NOR2xp5_ASAP7_6t_L U1008 ( .A(n92), .B(n301), .Y(n674) );
  XOR2xp5r_ASAP7_6t_L U1009 ( .A(n714), .B(n666), .Y(n704) );
  NAND2xp5R_ASAP7_6t_L U1010 ( .A(b[12]), .B(a[11]), .Y(n666) );
  NAND2xp5R_ASAP7_6t_L U1011 ( .A(b[13]), .B(a[10]), .Y(n714) );
  INVx1_ASAP7_6t_L U1012 ( .A(n698), .Y(n695) );
  XOR2xp5r_ASAP7_6t_L U1013 ( .A(n686), .B(n684), .Y(n689) );
  AO21x1_ASAP7_6t_L U1014 ( .A1(n715), .A2(n716), .B(n717), .Y(n684) );
  NOR3x1f_ASAP7_6t_L U1015 ( .A(n716), .B(n104), .C(n345), .Y(n717) );
  INVx1_ASAP7_6t_L U1016 ( .A(n685), .Y(n686) );
  XOR2xp5r_ASAP7_6t_L U1017 ( .A(n718), .B(n679), .Y(n685) );
  XOR2xp5r_ASAP7_6t_L U1018 ( .A(n678), .B(n719), .Y(n679) );
  NAND2xp5R_ASAP7_6t_L U1019 ( .A(b[10]), .B(a[13]), .Y(n719) );
  NOR2xp5_ASAP7_6t_L U1020 ( .A(n386), .B(n242), .Y(n678) );
  XOR2xp5r_ASAP7_6t_L U1021 ( .A(n720), .B(n687), .Y(n718) );
  NOR2xp5_ASAP7_6t_L U1022 ( .A(n345), .B(n91), .Y(n687) );
  NAND2xp5R_ASAP7_6t_L U1023 ( .A(b[9]), .B(a[14]), .Y(n720) );
  AOI22xp25_ASAP7_6t_L U1024 ( .A1(n721), .A2(n722), .B1(n723), .B2(n724), .Y(
        n693) );
  INVx1_ASAP7_6t_L U1025 ( .A(n722), .Y(n723) );
  AOI22xp25_ASAP7_6t_L U1026 ( .A1(n725), .A2(n726), .B1(n727), .B2(n728), .Y(
        n78) );
  INVx1_ASAP7_6t_L U1027 ( .A(n726), .Y(n727) );
  OAI22xp5_ASAP7_6t_L U1028 ( .A1(n79), .A2(n80), .B1(n729), .B2(n730), .Y(
        c[104]) );
  INVx1_ASAP7_6t_L U1029 ( .A(n729), .Y(n80) );
  XOR2xp5r_ASAP7_6t_L U1030 ( .A(n730), .B(n731), .Y(n729) );
  XOR2xp5r_ASAP7_6t_L U1031 ( .A(n728), .B(n726), .Y(n731) );
  AOI22xp25_ASAP7_6t_L U1032 ( .A1(n732), .A2(n733), .B1(n734), .B2(n735), .Y(
        n726) );
  XOR2xp5r_ASAP7_6t_L U1033 ( .A(n736), .B(n725), .Y(n734) );
  XOR2xp5r_ASAP7_6t_L U1034 ( .A(n737), .B(n725), .Y(n733) );
  XOR2xp5r_ASAP7_6t_L U1035 ( .A(n700), .B(n698), .Y(n725) );
  XOR2xp5r_ASAP7_6t_L U1036 ( .A(n738), .B(n702), .Y(n698) );
  AOI22xp25_ASAP7_6t_L U1037 ( .A1(n739), .A2(n740), .B1(n741), .B2(n742), .Y(
        n702) );
  XOR2xp5r_ASAP7_6t_L U1038 ( .A(n743), .B(n701), .Y(n742) );
  XOR2xp5r_ASAP7_6t_L U1039 ( .A(n744), .B(n701), .Y(n740) );
  XOR2xp5r_ASAP7_6t_L U1040 ( .A(n705), .B(n710), .Y(n701) );
  AO21x1_ASAP7_6t_L U1041 ( .A1(n745), .A2(n746), .B(n747), .Y(n710) );
  NOR3x1f_ASAP7_6t_L U1042 ( .A(n746), .B(n301), .C(n581), .Y(n747) );
  XOR2xp5r_ASAP7_6t_L U1043 ( .A(n748), .B(n712), .Y(n705) );
  XOR2xp5r_ASAP7_6t_L U1044 ( .A(n749), .B(n711), .Y(n712) );
  NOR2xp5_ASAP7_6t_L U1045 ( .A(n92), .B(n275), .Y(n711) );
  NAND2xp5R_ASAP7_6t_L U1046 ( .A(a[8]), .B(b[14]), .Y(n749) );
  XOR2xp5r_ASAP7_6t_L U1047 ( .A(n750), .B(n709), .Y(n748) );
  NOR2xp5_ASAP7_6t_L U1048 ( .A(n336), .B(n232), .Y(n709) );
  NAND2xp5R_ASAP7_6t_L U1049 ( .A(b[13]), .B(a[9]), .Y(n750) );
  XOR2xp5r_ASAP7_6t_L U1050 ( .A(n751), .B(n699), .Y(n738) );
  AOI22xp25_ASAP7_6t_L U1051 ( .A1(n752), .A2(n753), .B1(n754), .B2(n755), .Y(
        n699) );
  INVx1_ASAP7_6t_L U1052 ( .A(n756), .Y(n753) );
  NAND2xp5R_ASAP7_6t_L U1053 ( .A(b[11]), .B(a[11]), .Y(n751) );
  OA22x1_ASAP7_6t_L U1054 ( .A1(n757), .A2(n758), .B1(n759), .B2(n760), .Y(
        n700) );
  XOR2xp5r_ASAP7_6t_L U1055 ( .A(n722), .B(n721), .Y(n728) );
  AO21x1_ASAP7_6t_L U1056 ( .A1(n761), .A2(n762), .B(n763), .Y(n721) );
  NOR3x1f_ASAP7_6t_L U1057 ( .A(n762), .B(n104), .C(n212), .Y(n763) );
  XOR2xp5r_ASAP7_6t_L U1058 ( .A(n716), .B(n764), .Y(n722) );
  XOR2xp5r_ASAP7_6t_L U1059 ( .A(n724), .B(n765), .Y(n764) );
  NAND2xp5R_ASAP7_6t_L U1060 ( .A(b[8]), .B(a[14]), .Y(n765) );
  NOR2xp5_ASAP7_6t_L U1061 ( .A(n212), .B(n91), .Y(n724) );
  XOR2xp5r_ASAP7_6t_L U1062 ( .A(n715), .B(n766), .Y(n716) );
  NAND2xp5R_ASAP7_6t_L U1063 ( .A(b[9]), .B(a[13]), .Y(n766) );
  NOR2xp5_ASAP7_6t_L U1064 ( .A(n265), .B(n242), .Y(n715) );
  AOI22xp25_ASAP7_6t_L U1065 ( .A1(n767), .A2(n768), .B1(n769), .B2(n770), .Y(
        n730) );
  INVx1_ASAP7_6t_L U1066 ( .A(n768), .Y(n769) );
  AOI22xp25_ASAP7_6t_L U1067 ( .A1(n771), .A2(n772), .B1(n773), .B2(n774), .Y(
        n79) );
  OAI22xp5_ASAP7_6t_L U1068 ( .A1(n81), .A2(n82), .B1(n775), .B2(n776), .Y(
        c[103]) );
  INVx1_ASAP7_6t_L U1069 ( .A(n775), .Y(n82) );
  XOR2xp5r_ASAP7_6t_L U1070 ( .A(n776), .B(n777), .Y(n775) );
  XOR2xp5r_ASAP7_6t_L U1071 ( .A(n772), .B(n773), .Y(n777) );
  INVx1_ASAP7_6t_L U1072 ( .A(n771), .Y(n773) );
  OAI22xp5_ASAP7_6t_L U1073 ( .A1(n778), .A2(n779), .B1(n780), .B2(n781), .Y(
        n771) );
  XOR2xp5r_ASAP7_6t_L U1074 ( .A(n782), .B(n774), .Y(n781) );
  XOR2xp5r_ASAP7_6t_L U1075 ( .A(n783), .B(n774), .Y(n779) );
  XOR2xp5r_ASAP7_6t_L U1076 ( .A(n736), .B(n735), .Y(n774) );
  INVx1_ASAP7_6t_L U1077 ( .A(n732), .Y(n735) );
  XOR2xp5r_ASAP7_6t_L U1078 ( .A(n737), .B(n784), .Y(n732) );
  XOR2xp5r_ASAP7_6t_L U1079 ( .A(n758), .B(n759), .Y(n784) );
  INVx1_ASAP7_6t_L U1080 ( .A(n757), .Y(n759) );
  AOI22xp25_ASAP7_6t_L U1081 ( .A1(n785), .A2(n786), .B1(n787), .B2(n788), .Y(
        n757) );
  XOR2xp5r_ASAP7_6t_L U1082 ( .A(n789), .B(n760), .Y(n788) );
  XOR2xp5r_ASAP7_6t_L U1083 ( .A(n790), .B(n760), .Y(n786) );
  XOR2xp5r_ASAP7_6t_L U1084 ( .A(n741), .B(n744), .Y(n760) );
  AO21x1_ASAP7_6t_L U1085 ( .A1(n791), .A2(n792), .B(n793), .Y(n744) );
  NOR3x1f_ASAP7_6t_L U1086 ( .A(n792), .B(n275), .C(n581), .Y(n793) );
  INVx1_ASAP7_6t_L U1087 ( .A(n739), .Y(n741) );
  XOR2xp5r_ASAP7_6t_L U1088 ( .A(n794), .B(n746), .Y(n739) );
  XOR2xp5r_ASAP7_6t_L U1089 ( .A(n795), .B(n745), .Y(n746) );
  NOR2xp5_ASAP7_6t_L U1090 ( .A(n92), .B(n213), .Y(n745) );
  NAND2xp5R_ASAP7_6t_L U1091 ( .A(a[7]), .B(b[14]), .Y(n795) );
  XOR2xp5r_ASAP7_6t_L U1092 ( .A(n796), .B(n743), .Y(n794) );
  NOR2xp5_ASAP7_6t_L U1093 ( .A(n336), .B(n356), .Y(n743) );
  NAND2xp5R_ASAP7_6t_L U1094 ( .A(b[13]), .B(a[8]), .Y(n796) );
  XOR2xp5r_ASAP7_6t_L U1095 ( .A(n752), .B(n756), .Y(n758) );
  AOI21xp25_ASAP7_6t_L U1096 ( .A1(n797), .A2(n798), .B(n799), .Y(n756) );
  NOR3x1f_ASAP7_6t_L U1097 ( .A(n798), .B(n236), .C(n277), .Y(n799) );
  XOR2xp5r_ASAP7_6t_L U1098 ( .A(n755), .B(n754), .Y(n752) );
  NOR2xp5_ASAP7_6t_L U1099 ( .A(n386), .B(n232), .Y(n754) );
  NOR2xp5_ASAP7_6t_L U1100 ( .A(n265), .B(n236), .Y(n755) );
  AO22x1_ASAP7_6t_L U1101 ( .A1(n800), .A2(n801), .B1(n802), .B2(n803), .Y(
        n737) );
  INVx1_ASAP7_6t_L U1102 ( .A(n802), .Y(n801) );
  OAI22xp5_ASAP7_6t_L U1103 ( .A1(n804), .A2(n805), .B1(n806), .B2(n807), .Y(
        n736) );
  XOR2xp5r_ASAP7_6t_L U1104 ( .A(n767), .B(n768), .Y(n772) );
  XOR2xp5r_ASAP7_6t_L U1105 ( .A(n762), .B(n808), .Y(n768) );
  XOR2xp5r_ASAP7_6t_L U1106 ( .A(n770), .B(n809), .Y(n808) );
  NAND2xp5R_ASAP7_6t_L U1107 ( .A(b[7]), .B(a[14]), .Y(n809) );
  NOR2xp5_ASAP7_6t_L U1108 ( .A(n272), .B(n91), .Y(n770) );
  XOR2xp5r_ASAP7_6t_L U1109 ( .A(n810), .B(n761), .Y(n762) );
  NOR2xp5_ASAP7_6t_L U1110 ( .A(n277), .B(n242), .Y(n761) );
  NAND2xp5R_ASAP7_6t_L U1111 ( .A(a[13]), .B(b[8]), .Y(n810) );
  OR2x2_ASAP7_6t_L U1112 ( .A(n811), .B(n812), .Y(n767) );
  NOR3x1f_ASAP7_6t_L U1113 ( .A(n813), .B(n102), .C(n212), .Y(n812) );
  NOR3x1f_ASAP7_6t_L U1114 ( .A(n814), .B(n104), .C(n272), .Y(n811) );
  OA22x1_ASAP7_6t_L U1115 ( .A1(n815), .A2(n816), .B1(n817), .B2(n818), .Y(
        n776) );
  INVx1_ASAP7_6t_L U1116 ( .A(n817), .Y(n815) );
  AOI22xp25_ASAP7_6t_L U1117 ( .A1(n819), .A2(n820), .B1(n821), .B2(n822), .Y(
        n81) );
  INVx1_ASAP7_6t_L U1118 ( .A(n822), .Y(n819) );
  OAI22xp5_ASAP7_6t_L U1119 ( .A1(n823), .A2(n824), .B1(n84), .B2(n83), .Y(
        c[102]) );
  AOI22xp25_ASAP7_6t_L U1120 ( .A1(n825), .A2(n826), .B1(n827), .B2(n828), .Y(
        n83) );
  INVx1_ASAP7_6t_L U1121 ( .A(n825), .Y(n827) );
  INVx1_ASAP7_6t_L U1122 ( .A(n84), .Y(n824) );
  XOR2xp5r_ASAP7_6t_L U1123 ( .A(n823), .B(n829), .Y(n84) );
  XOR2xp5r_ASAP7_6t_L U1124 ( .A(n821), .B(n822), .Y(n829) );
  OAI22xp5_ASAP7_6t_L U1125 ( .A1(n830), .A2(n831), .B1(n832), .B2(n833), .Y(
        n822) );
  XOR2xp5r_ASAP7_6t_L U1126 ( .A(n834), .B(n820), .Y(n833) );
  XOR2xp5r_ASAP7_6t_L U1127 ( .A(n835), .B(n820), .Y(n831) );
  XOR2xp5r_ASAP7_6t_L U1128 ( .A(n783), .B(n778), .Y(n820) );
  INVx1_ASAP7_6t_L U1129 ( .A(n780), .Y(n778) );
  XOR2xp5r_ASAP7_6t_L U1130 ( .A(n782), .B(n836), .Y(n780) );
  XOR2xp5r_ASAP7_6t_L U1131 ( .A(n805), .B(n806), .Y(n836) );
  INVx1_ASAP7_6t_L U1132 ( .A(n804), .Y(n806) );
  AOI22xp25_ASAP7_6t_L U1133 ( .A1(n837), .A2(n838), .B1(n839), .B2(n840), .Y(
        n804) );
  XOR2xp5r_ASAP7_6t_L U1134 ( .A(n841), .B(n807), .Y(n840) );
  XOR2xp5r_ASAP7_6t_L U1135 ( .A(n842), .B(n807), .Y(n838) );
  XOR2xp5r_ASAP7_6t_L U1136 ( .A(n785), .B(n790), .Y(n807) );
  AOI21xp25_ASAP7_6t_L U1137 ( .A1(n843), .A2(n844), .B(n845), .Y(n790) );
  NOR3x1f_ASAP7_6t_L U1138 ( .A(n844), .B(n213), .C(n581), .Y(n845) );
  INVx1_ASAP7_6t_L U1139 ( .A(n787), .Y(n785) );
  XOR2xp5r_ASAP7_6t_L U1140 ( .A(n792), .B(n846), .Y(n787) );
  XOR2xp5r_ASAP7_6t_L U1141 ( .A(n789), .B(n847), .Y(n846) );
  NAND2xp5R_ASAP7_6t_L U1142 ( .A(b[13]), .B(a[7]), .Y(n847) );
  NAND2xp5R_ASAP7_6t_L U1143 ( .A(b[12]), .B(a[8]), .Y(n789) );
  XOR2xp5r_ASAP7_6t_L U1144 ( .A(n791), .B(n848), .Y(n792) );
  NAND2xp5R_ASAP7_6t_L U1145 ( .A(b[14]), .B(a[6]), .Y(n848) );
  NOR2xp5_ASAP7_6t_L U1146 ( .A(n92), .B(n390), .Y(n791) );
  XOR2xp5r_ASAP7_6t_L U1147 ( .A(n802), .B(n800), .Y(n805) );
  AO21x1_ASAP7_6t_L U1148 ( .A1(n849), .A2(n850), .B(n851), .Y(n800) );
  NOR3x1f_ASAP7_6t_L U1149 ( .A(n850), .B(n232), .C(n277), .Y(n851) );
  XOR2xp5r_ASAP7_6t_L U1150 ( .A(n798), .B(n852), .Y(n802) );
  XOR2xp5r_ASAP7_6t_L U1151 ( .A(n853), .B(n803), .Y(n852) );
  NOR2xp5_ASAP7_6t_L U1152 ( .A(n345), .B(n242), .Y(n803) );
  NOR2xp5_ASAP7_6t_L U1153 ( .A(n236), .B(n277), .Y(n853) );
  XOR2xp5r_ASAP7_6t_L U1154 ( .A(n854), .B(n797), .Y(n798) );
  NOR2xp5_ASAP7_6t_L U1155 ( .A(n386), .B(n356), .Y(n797) );
  NAND2xp5R_ASAP7_6t_L U1156 ( .A(a[10]), .B(b[10]), .Y(n854) );
  AOI22xp25_ASAP7_6t_L U1157 ( .A1(n855), .A2(n856), .B1(n857), .B2(n858), .Y(
        n782) );
  OA22x1_ASAP7_6t_L U1158 ( .A1(n859), .A2(n860), .B1(n861), .B2(n862), .Y(
        n783) );
  INVx1_ASAP7_6t_L U1159 ( .A(n861), .Y(n859) );
  XOR2xp5r_ASAP7_6t_L U1160 ( .A(n817), .B(n818), .Y(n821) );
  AOI21xp25_ASAP7_6t_L U1161 ( .A1(n863), .A2(n864), .B(n865), .Y(n818) );
  NOR3x1f_ASAP7_6t_L U1162 ( .A(n864), .B(n104), .C(n302), .Y(n865) );
  XOR2xp5r_ASAP7_6t_L U1163 ( .A(n866), .B(n814), .Y(n817) );
  INVx1_ASAP7_6t_L U1164 ( .A(n813), .Y(n814) );
  XOR2xp5r_ASAP7_6t_L U1165 ( .A(n867), .B(n868), .Y(n813) );
  NAND2xp5R_ASAP7_6t_L U1166 ( .A(b[7]), .B(a[13]), .Y(n868) );
  AOI22xp25_ASAP7_6t_L U1167 ( .A1(n869), .A2(n870), .B1(n871), .B2(n872), .Y(
        n867) );
  XOR2xp5r_ASAP7_6t_L U1168 ( .A(n873), .B(n816), .Y(n866) );
  NAND2xp5R_ASAP7_6t_L U1169 ( .A(b[5]), .B(a[15]), .Y(n816) );
  NAND2xp5R_ASAP7_6t_L U1170 ( .A(b[6]), .B(a[14]), .Y(n873) );
  OA22x1_ASAP7_6t_L U1171 ( .A1(n874), .A2(n875), .B1(n876), .B2(n877), .Y(
        n823) );
  INVx1_ASAP7_6t_L U1172 ( .A(n875), .Y(n876) );
  OAI22xp5_ASAP7_6t_L U1173 ( .A1(n85), .A2(n86), .B1(n878), .B2(n879), .Y(
        c[101]) );
  INVx1_ASAP7_6t_L U1174 ( .A(n86), .Y(n878) );
  XOR2xp5r_ASAP7_6t_L U1175 ( .A(n879), .B(n880), .Y(n86) );
  XOR2xp5r_ASAP7_6t_L U1176 ( .A(n826), .B(n825), .Y(n880) );
  OAI22xp5_ASAP7_6t_L U1177 ( .A1(n881), .A2(n882), .B1(n883), .B2(n884), .Y(
        n825) );
  XOR2xp5r_ASAP7_6t_L U1178 ( .A(n885), .B(n828), .Y(n884) );
  INVx1_ASAP7_6t_L U1179 ( .A(n881), .Y(n883) );
  XOR2xp5r_ASAP7_6t_L U1180 ( .A(n886), .B(n828), .Y(n882) );
  XOR2xp5r_ASAP7_6t_L U1181 ( .A(n835), .B(n830), .Y(n828) );
  INVx1_ASAP7_6t_L U1182 ( .A(n832), .Y(n830) );
  XOR2xp5r_ASAP7_6t_L U1183 ( .A(n834), .B(n887), .Y(n832) );
  XOR2xp5r_ASAP7_6t_L U1184 ( .A(n860), .B(n861), .Y(n887) );
  OAI22xp5_ASAP7_6t_L U1185 ( .A1(n888), .A2(n889), .B1(n890), .B2(n891), .Y(
        n861) );
  XOR2xp5r_ASAP7_6t_L U1186 ( .A(n892), .B(n862), .Y(n891) );
  XOR2xp5r_ASAP7_6t_L U1187 ( .A(n893), .B(n862), .Y(n889) );
  XOR2xp5r_ASAP7_6t_L U1188 ( .A(n837), .B(n842), .Y(n862) );
  AOI21xp25_ASAP7_6t_L U1189 ( .A1(n894), .A2(n895), .B(n896), .Y(n842) );
  NOR3x1f_ASAP7_6t_L U1190 ( .A(n895), .B(n390), .C(n581), .Y(n896) );
  INVx1_ASAP7_6t_L U1191 ( .A(n839), .Y(n837) );
  XOR2xp5r_ASAP7_6t_L U1192 ( .A(n897), .B(n844), .Y(n839) );
  XOR2xp5r_ASAP7_6t_L U1193 ( .A(n898), .B(n843), .Y(n844) );
  NOR2xp5_ASAP7_6t_L U1194 ( .A(n92), .B(n278), .Y(n843) );
  NAND2xp5R_ASAP7_6t_L U1195 ( .A(a[5]), .B(b[14]), .Y(n898) );
  XOR2xp5r_ASAP7_6t_L U1196 ( .A(n899), .B(n841), .Y(n897) );
  NAND2xp5R_ASAP7_6t_L U1197 ( .A(b[12]), .B(a[7]), .Y(n841) );
  NAND2xp5R_ASAP7_6t_L U1198 ( .A(b[13]), .B(a[6]), .Y(n899) );
  XOR2xp5r_ASAP7_6t_L U1199 ( .A(n857), .B(n855), .Y(n860) );
  AO21x1_ASAP7_6t_L U1200 ( .A1(n900), .A2(n901), .B(n902), .Y(n855) );
  NOR3x1f_ASAP7_6t_L U1201 ( .A(n901), .B(n356), .C(n277), .Y(n902) );
  INVx1_ASAP7_6t_L U1202 ( .A(n856), .Y(n857) );
  XOR2xp5r_ASAP7_6t_L U1203 ( .A(n903), .B(n850), .Y(n856) );
  XOR2xp5r_ASAP7_6t_L U1204 ( .A(n904), .B(n849), .Y(n850) );
  NOR2xp5_ASAP7_6t_L U1205 ( .A(n386), .B(n301), .Y(n849) );
  NAND2xp5R_ASAP7_6t_L U1206 ( .A(a[9]), .B(b[10]), .Y(n904) );
  XOR2xp5r_ASAP7_6t_L U1207 ( .A(n905), .B(n858), .Y(n903) );
  NOR2xp5_ASAP7_6t_L U1208 ( .A(n345), .B(n236), .Y(n858) );
  NAND2xp5R_ASAP7_6t_L U1209 ( .A(b[9]), .B(a[10]), .Y(n905) );
  AOI22xp25_ASAP7_6t_L U1210 ( .A1(n906), .A2(n907), .B1(n908), .B2(n909), .Y(
        n834) );
  INVx1_ASAP7_6t_L U1211 ( .A(n908), .Y(n907) );
  OA22x1_ASAP7_6t_L U1212 ( .A1(n910), .A2(n911), .B1(n912), .B2(n913), .Y(
        n835) );
  XOR2xp5r_ASAP7_6t_L U1213 ( .A(n874), .B(n875), .Y(n826) );
  XOR2xp5r_ASAP7_6t_L U1214 ( .A(n914), .B(n864), .Y(n875) );
  OA22x1_ASAP7_6t_L U1215 ( .A1(n915), .A2(n916), .B1(n917), .B2(n918), .Y(
        n864) );
  XOR2xp5r_ASAP7_6t_L U1216 ( .A(n919), .B(n920), .Y(n918) );
  XOR2xp5r_ASAP7_6t_L U1217 ( .A(n921), .B(n920), .Y(n916) );
  INVx1_ASAP7_6t_L U1218 ( .A(n863), .Y(n920) );
  XOR2xp5r_ASAP7_6t_L U1219 ( .A(n872), .B(n871), .Y(n863) );
  AO21x1_ASAP7_6t_L U1220 ( .A1(n922), .A2(n923), .B(n924), .Y(n871) );
  NOR3x1f_ASAP7_6t_L U1221 ( .A(n923), .B(n102), .C(n302), .Y(n924) );
  INVx1_ASAP7_6t_L U1222 ( .A(b[5]), .Y(n302) );
  XOR2xp5r_ASAP7_6t_L U1223 ( .A(n870), .B(n869), .Y(n872) );
  NOR2xp5_ASAP7_6t_L U1224 ( .A(n272), .B(n102), .Y(n869) );
  NOR2xp5_ASAP7_6t_L U1225 ( .A(n212), .B(n242), .Y(n870) );
  INVx1_ASAP7_6t_L U1226 ( .A(n917), .Y(n915) );
  XOR2xp5r_ASAP7_6t_L U1227 ( .A(n925), .B(n877), .Y(n914) );
  NAND2xp5R_ASAP7_6t_L U1228 ( .A(b[4]), .B(a[15]), .Y(n877) );
  NAND2xp5R_ASAP7_6t_L U1229 ( .A(b[5]), .B(a[14]), .Y(n925) );
  AOI21xp25_ASAP7_6t_L U1230 ( .A1(n926), .A2(n927), .B(n928), .Y(n874) );
  NOR3x1f_ASAP7_6t_L U1231 ( .A(n927), .B(n231), .C(n91), .Y(n928) );
  AOI22xp25_ASAP7_6t_L U1232 ( .A1(n929), .A2(n930), .B1(n931), .B2(n932), .Y(
        n879) );
  AOI22xp25_ASAP7_6t_L U1233 ( .A1(n933), .A2(n934), .B1(n935), .B2(n936), .Y(
        n85) );
  INVx1_ASAP7_6t_L U1234 ( .A(n936), .Y(n933) );
  OAI22xp5_ASAP7_6t_L U1235 ( .A1(n937), .A2(n938), .B1(n88), .B2(n87), .Y(
        c[100]) );
  AOI22xp25_ASAP7_6t_L U1236 ( .A1(n114), .A2(n939), .B1(n115), .B2(n940), .Y(
        n87) );
  XOR2xp5r_ASAP7_6t_L U1237 ( .A(n941), .B(n942), .Y(n115) );
  INVx1_ASAP7_6t_L U1238 ( .A(n940), .Y(n114) );
  OAI22xp5_ASAP7_6t_L U1239 ( .A1(n943), .A2(n944), .B1(n130), .B2(n945), .Y(
        n940) );
  XOR2xp5r_ASAP7_6t_L U1240 ( .A(n946), .B(n939), .Y(n945) );
  INVx1_ASAP7_6t_L U1241 ( .A(n943), .Y(n130) );
  XOR2xp5r_ASAP7_6t_L U1242 ( .A(n129), .B(n939), .Y(n944) );
  XOR2xp5r_ASAP7_6t_L U1243 ( .A(n947), .B(n948), .Y(n939) );
  AOI22xp25_ASAP7_6t_L U1244 ( .A1(n949), .A2(n157), .B1(n156), .B2(n950), .Y(
        n129) );
  XOR2xp5r_ASAP7_6t_L U1245 ( .A(n951), .B(n952), .Y(n157) );
  INVx1_ASAP7_6t_L U1246 ( .A(n156), .Y(n949) );
  AOI22xp25_ASAP7_6t_L U1247 ( .A1(n953), .A2(n954), .B1(n207), .B2(n955), .Y(
        n156) );
  XOR2xp5r_ASAP7_6t_L U1248 ( .A(n956), .B(n950), .Y(n955) );
  INVx1_ASAP7_6t_L U1249 ( .A(n953), .Y(n207) );
  XOR2xp5r_ASAP7_6t_L U1250 ( .A(n208), .B(n950), .Y(n954) );
  XOR2xp5r_ASAP7_6t_L U1251 ( .A(n957), .B(n958), .Y(n950) );
  AO21x1_ASAP7_6t_L U1252 ( .A1(n959), .A2(n266), .B(n960), .Y(n208) );
  NOR3x1f_ASAP7_6t_L U1253 ( .A(n266), .B(n386), .C(n90), .Y(n960) );
  XOR2xp5r_ASAP7_6t_L U1254 ( .A(n961), .B(n959), .Y(n266) );
  NAND2xp5R_ASAP7_6t_L U1255 ( .A(a[1]), .B(b[12]), .Y(n961) );
  NOR2xp5_ASAP7_6t_L U1256 ( .A(n94), .B(n581), .Y(n959) );
  INVx1_ASAP7_6t_L U1257 ( .A(b[13]), .Y(n581) );
  XOR2xp5r_ASAP7_6t_L U1258 ( .A(n962), .B(n963), .Y(n953) );
  XOR2xp5r_ASAP7_6t_L U1259 ( .A(n956), .B(n964), .Y(n963) );
  NAND2xp5R_ASAP7_6t_L U1260 ( .A(b[12]), .B(a[2]), .Y(n964) );
  NOR2xp5_ASAP7_6t_L U1261 ( .A(n428), .B(n386), .Y(n956) );
  XOR2xp5r_ASAP7_6t_L U1262 ( .A(n946), .B(n965), .Y(n943) );
  XOR2xp5r_ASAP7_6t_L U1263 ( .A(n966), .B(n967), .Y(n965) );
  AOI21xp25_ASAP7_6t_L U1264 ( .A1(n951), .A2(n952), .B(n968), .Y(n946) );
  NOR3x1f_ASAP7_6t_L U1265 ( .A(n951), .B(n345), .C(n275), .Y(n968) );
  AO21x1_ASAP7_6t_L U1266 ( .A1(n969), .A2(n215), .B(n970), .Y(n952) );
  NOR3x1f_ASAP7_6t_L U1267 ( .A(n215), .B(n213), .C(n345), .Y(n970) );
  XOR2xp5r_ASAP7_6t_L U1268 ( .A(n971), .B(n969), .Y(n215) );
  NAND2xp5R_ASAP7_6t_L U1269 ( .A(a[5]), .B(b[9]), .Y(n971) );
  NOR2xp5_ASAP7_6t_L U1270 ( .A(n265), .B(n278), .Y(n969) );
  XOR2xp5r_ASAP7_6t_L U1271 ( .A(n972), .B(n973), .Y(n951) );
  XOR2xp5r_ASAP7_6t_L U1272 ( .A(n974), .B(n975), .Y(n973) );
  NOR2xp5_ASAP7_6t_L U1273 ( .A(n345), .B(n275), .Y(n974) );
  INVx1_ASAP7_6t_L U1274 ( .A(n88), .Y(n938) );
  XOR2xp5r_ASAP7_6t_L U1275 ( .A(n937), .B(n976), .Y(n88) );
  XOR2xp5r_ASAP7_6t_L U1276 ( .A(n935), .B(n936), .Y(n976) );
  OAI22xp5_ASAP7_6t_L U1277 ( .A1(n947), .A2(n977), .B1(n978), .B2(n979), .Y(
        n936) );
  XOR2xp5r_ASAP7_6t_L U1278 ( .A(n980), .B(n934), .Y(n979) );
  INVx1_ASAP7_6t_L U1279 ( .A(n947), .Y(n978) );
  XOR2xp5r_ASAP7_6t_L U1280 ( .A(n948), .B(n934), .Y(n977) );
  XOR2xp5r_ASAP7_6t_L U1281 ( .A(n886), .B(n881), .Y(n934) );
  XOR2xp5r_ASAP7_6t_L U1282 ( .A(n885), .B(n981), .Y(n881) );
  XOR2xp5r_ASAP7_6t_L U1283 ( .A(n911), .B(n910), .Y(n981) );
  INVx1_ASAP7_6t_L U1284 ( .A(n912), .Y(n910) );
  XOR2xp5r_ASAP7_6t_L U1285 ( .A(n982), .B(n913), .Y(n912) );
  XOR2xp5r_ASAP7_6t_L U1286 ( .A(n888), .B(n893), .Y(n913) );
  OAI22xp5_ASAP7_6t_L U1287 ( .A1(n983), .A2(n984), .B1(n985), .B2(n986), .Y(
        n893) );
  INVx1_ASAP7_6t_L U1288 ( .A(n983), .Y(n985) );
  INVx1_ASAP7_6t_L U1289 ( .A(n890), .Y(n888) );
  XOR2xp5r_ASAP7_6t_L U1290 ( .A(n987), .B(n895), .Y(n890) );
  XOR2xp5r_ASAP7_6t_L U1291 ( .A(n988), .B(n894), .Y(n895) );
  NOR2xp5_ASAP7_6t_L U1292 ( .A(n428), .B(n92), .Y(n894) );
  INVx1_ASAP7_6t_L U1293 ( .A(b[15]), .Y(n92) );
  NAND2xp5R_ASAP7_6t_L U1294 ( .A(a[4]), .B(b[14]), .Y(n988) );
  XOR2xp5r_ASAP7_6t_L U1295 ( .A(n989), .B(n892), .Y(n987) );
  NOR2xp5_ASAP7_6t_L U1296 ( .A(n336), .B(n213), .Y(n892) );
  NAND2xp5R_ASAP7_6t_L U1297 ( .A(b[13]), .B(a[5]), .Y(n989) );
  AOI21xp25_ASAP7_6t_L U1298 ( .A1(n990), .A2(n991), .B(n992), .Y(n982) );
  NOR3x1f_ASAP7_6t_L U1299 ( .A(n990), .B(n390), .C(n336), .Y(n992) );
  XOR2xp5r_ASAP7_6t_L U1300 ( .A(n908), .B(n906), .Y(n911) );
  OAI22xp5_ASAP7_6t_L U1301 ( .A1(n993), .A2(n994), .B1(n995), .B2(n996), .Y(
        n906) );
  XOR2xp5r_ASAP7_6t_L U1302 ( .A(n901), .B(n997), .Y(n908) );
  XOR2xp5r_ASAP7_6t_L U1303 ( .A(n998), .B(n909), .Y(n997) );
  NOR2xp5_ASAP7_6t_L U1304 ( .A(n345), .B(n232), .Y(n909) );
  NOR2xp5_ASAP7_6t_L U1305 ( .A(n356), .B(n277), .Y(n998) );
  INVx1_ASAP7_6t_L U1306 ( .A(b[9]), .Y(n277) );
  XOR2xp5r_ASAP7_6t_L U1307 ( .A(n999), .B(n900), .Y(n901) );
  NOR2xp5_ASAP7_6t_L U1308 ( .A(n275), .B(n386), .Y(n900) );
  INVx1_ASAP7_6t_L U1309 ( .A(b[11]), .Y(n386) );
  NAND2xp5R_ASAP7_6t_L U1310 ( .A(a[8]), .B(b[10]), .Y(n999) );
  AOI21xp25_ASAP7_6t_L U1311 ( .A1(n1000), .A2(n1001), .B(n1002), .Y(n885) );
  NOR3x1f_ASAP7_6t_L U1312 ( .A(n1000), .B(n356), .C(n345), .Y(n1002) );
  AOI22xp25_ASAP7_6t_L U1313 ( .A1(n1003), .A2(n1004), .B1(n1005), .B2(n1006), 
        .Y(n886) );
  AOI22xp25_ASAP7_6t_L U1314 ( .A1(n967), .A2(n966), .B1(n1007), .B2(n1008), 
        .Y(n948) );
  XOR2xp5r_ASAP7_6t_L U1315 ( .A(n1009), .B(n1010), .Y(n966) );
  INVx1_ASAP7_6t_L U1316 ( .A(n1007), .Y(n967) );
  XOR2xp5r_ASAP7_6t_L U1317 ( .A(n1011), .B(n1008), .Y(n1007) );
  XOR2xp5r_ASAP7_6t_L U1318 ( .A(n1012), .B(n1013), .Y(n1008) );
  AOI21xp25_ASAP7_6t_L U1319 ( .A1(n957), .A2(n958), .B(n1014), .Y(n1011) );
  NOR3x1f_ASAP7_6t_L U1320 ( .A(n957), .B(n336), .C(n428), .Y(n1014) );
  AO21x1_ASAP7_6t_L U1321 ( .A1(n1015), .A2(n962), .B(n1016), .Y(n958) );
  NOR3x1f_ASAP7_6t_L U1322 ( .A(n962), .B(n90), .C(n336), .Y(n1016) );
  INVx1_ASAP7_6t_L U1323 ( .A(a[2]), .Y(n90) );
  XOR2xp5r_ASAP7_6t_L U1324 ( .A(n1015), .B(n1017), .Y(n962) );
  NAND2xp5R_ASAP7_6t_L U1325 ( .A(b[13]), .B(a[1]), .Y(n1017) );
  NOR2xp5_ASAP7_6t_L U1326 ( .A(n98), .B(n94), .Y(n1015) );
  INVx1_ASAP7_6t_L U1327 ( .A(a[0]), .Y(n94) );
  XOR2xp5r_ASAP7_6t_L U1328 ( .A(n1018), .B(n1019), .Y(n957) );
  XOR2xp5r_ASAP7_6t_L U1329 ( .A(n1020), .B(n1021), .Y(n1019) );
  NOR2xp5_ASAP7_6t_L U1330 ( .A(n336), .B(n428), .Y(n1020) );
  XOR2xp5r_ASAP7_6t_L U1331 ( .A(n980), .B(n1022), .Y(n947) );
  XOR2xp5r_ASAP7_6t_L U1332 ( .A(n1004), .B(n1003), .Y(n1022) );
  INVx1_ASAP7_6t_L U1333 ( .A(n1005), .Y(n1003) );
  XOR2xp5r_ASAP7_6t_L U1334 ( .A(n1023), .B(n1006), .Y(n1005) );
  XOR2xp5r_ASAP7_6t_L U1335 ( .A(n990), .B(n991), .Y(n1006) );
  OAI22xp5_ASAP7_6t_L U1336 ( .A1(n1024), .A2(n1025), .B1(n1026), .B2(n1027), 
        .Y(n991) );
  XOR2xp5r_ASAP7_6t_L U1337 ( .A(n983), .B(n1028), .Y(n990) );
  XOR2xp5r_ASAP7_6t_L U1338 ( .A(n1029), .B(n984), .Y(n1028) );
  NAND2xp5R_ASAP7_6t_L U1339 ( .A(b[13]), .B(a[4]), .Y(n984) );
  NOR2xp5_ASAP7_6t_L U1340 ( .A(n390), .B(n336), .Y(n1029) );
  XOR2xp5r_ASAP7_6t_L U1341 ( .A(n1030), .B(n986), .Y(n983) );
  NAND2xp5R_ASAP7_6t_L U1342 ( .A(b[15]), .B(a[2]), .Y(n986) );
  NOR2xp5_ASAP7_6t_L U1343 ( .A(n98), .B(n428), .Y(n1030) );
  INVx1_ASAP7_6t_L U1344 ( .A(a[3]), .Y(n428) );
  AOI21xp25_ASAP7_6t_L U1345 ( .A1(n1012), .A2(n1013), .B(n1031), .Y(n1023) );
  NOR3x1f_ASAP7_6t_L U1346 ( .A(n1012), .B(n278), .C(n336), .Y(n1031) );
  OAI22xp5_ASAP7_6t_L U1347 ( .A1(n1018), .A2(n1021), .B1(n1032), .B2(n1033), 
        .Y(n1013) );
  INVx1_ASAP7_6t_L U1348 ( .A(n1018), .Y(n1032) );
  NAND2xp5R_ASAP7_6t_L U1349 ( .A(a[2]), .B(b[13]), .Y(n1021) );
  XOR2xp5r_ASAP7_6t_L U1350 ( .A(n1034), .B(n1033), .Y(n1018) );
  NAND2xp5R_ASAP7_6t_L U1351 ( .A(b[15]), .B(a[0]), .Y(n1033) );
  NOR2xp5_ASAP7_6t_L U1352 ( .A(n95), .B(n98), .Y(n1034) );
  INVx1_ASAP7_6t_L U1353 ( .A(b[14]), .Y(n98) );
  INVx1_ASAP7_6t_L U1354 ( .A(a[1]), .Y(n95) );
  XOR2xp5r_ASAP7_6t_L U1355 ( .A(n1024), .B(n1035), .Y(n1012) );
  XOR2xp5r_ASAP7_6t_L U1356 ( .A(n1036), .B(n1025), .Y(n1035) );
  NAND2xp5R_ASAP7_6t_L U1357 ( .A(a[3]), .B(b[13]), .Y(n1025) );
  NOR2xp5_ASAP7_6t_L U1358 ( .A(n278), .B(n336), .Y(n1036) );
  INVx1_ASAP7_6t_L U1359 ( .A(b[12]), .Y(n336) );
  INVx1_ASAP7_6t_L U1360 ( .A(a[4]), .Y(n278) );
  INVx1_ASAP7_6t_L U1361 ( .A(n1026), .Y(n1024) );
  XOR2xp5r_ASAP7_6t_L U1362 ( .A(n1027), .B(n1037), .Y(n1026) );
  NAND2xp5R_ASAP7_6t_L U1363 ( .A(a[2]), .B(b[14]), .Y(n1037) );
  NAND2xp5R_ASAP7_6t_L U1364 ( .A(b[15]), .B(a[1]), .Y(n1027) );
  XOR2xp5r_ASAP7_6t_L U1365 ( .A(n1000), .B(n1001), .Y(n1004) );
  OAI22xp5_ASAP7_6t_L U1366 ( .A1(n1038), .A2(n1039), .B1(n1040), .B2(n1041), 
        .Y(n1001) );
  INVx1_ASAP7_6t_L U1367 ( .A(n1038), .Y(n1040) );
  XOR2xp5r_ASAP7_6t_L U1368 ( .A(n1042), .B(n995), .Y(n1000) );
  INVx1_ASAP7_6t_L U1369 ( .A(n993), .Y(n995) );
  XOR2xp5r_ASAP7_6t_L U1370 ( .A(n1043), .B(n996), .Y(n993) );
  NAND2xp5R_ASAP7_6t_L U1371 ( .A(b[11]), .B(a[6]), .Y(n996) );
  NOR2xp5_ASAP7_6t_L U1372 ( .A(n265), .B(n275), .Y(n1043) );
  INVx1_ASAP7_6t_L U1373 ( .A(a[7]), .Y(n275) );
  XOR2xp5r_ASAP7_6t_L U1374 ( .A(n1044), .B(n994), .Y(n1042) );
  NAND2xp5R_ASAP7_6t_L U1375 ( .A(b[9]), .B(a[8]), .Y(n994) );
  NAND2xp5R_ASAP7_6t_L U1376 ( .A(b[8]), .B(a[9]), .Y(n1044) );
  AOI21xp25_ASAP7_6t_L U1377 ( .A1(n1009), .A2(n1010), .B(n1045), .Y(n980) );
  NOR3x1f_ASAP7_6t_L U1378 ( .A(n1009), .B(n301), .C(n345), .Y(n1045) );
  OAI22xp5_ASAP7_6t_L U1379 ( .A1(n972), .A2(n975), .B1(n1046), .B2(n1047), 
        .Y(n1010) );
  INVx1_ASAP7_6t_L U1380 ( .A(n972), .Y(n1046) );
  NAND2xp5R_ASAP7_6t_L U1381 ( .A(a[6]), .B(b[9]), .Y(n975) );
  XOR2xp5r_ASAP7_6t_L U1382 ( .A(n1048), .B(n1047), .Y(n972) );
  NAND2xp5R_ASAP7_6t_L U1383 ( .A(b[11]), .B(a[4]), .Y(n1047) );
  NOR2xp5_ASAP7_6t_L U1384 ( .A(n265), .B(n390), .Y(n1048) );
  INVx1_ASAP7_6t_L U1385 ( .A(a[5]), .Y(n390) );
  XOR2xp5r_ASAP7_6t_L U1386 ( .A(n1038), .B(n1049), .Y(n1009) );
  XOR2xp5r_ASAP7_6t_L U1387 ( .A(n1050), .B(n1039), .Y(n1049) );
  NAND2xp5R_ASAP7_6t_L U1388 ( .A(a[7]), .B(b[9]), .Y(n1039) );
  NOR2xp5_ASAP7_6t_L U1389 ( .A(n301), .B(n345), .Y(n1050) );
  INVx1_ASAP7_6t_L U1390 ( .A(b[8]), .Y(n345) );
  XOR2xp5r_ASAP7_6t_L U1391 ( .A(n1051), .B(n1041), .Y(n1038) );
  NAND2xp5R_ASAP7_6t_L U1392 ( .A(b[11]), .B(a[5]), .Y(n1041) );
  NOR2xp5_ASAP7_6t_L U1393 ( .A(n265), .B(n213), .Y(n1051) );
  INVx1_ASAP7_6t_L U1394 ( .A(a[6]), .Y(n213) );
  INVx1_ASAP7_6t_L U1395 ( .A(b[10]), .Y(n265) );
  XOR2xp5r_ASAP7_6t_L U1396 ( .A(n930), .B(n929), .Y(n935) );
  INVx1_ASAP7_6t_L U1397 ( .A(n932), .Y(n929) );
  XOR2xp5r_ASAP7_6t_L U1398 ( .A(n927), .B(n1052), .Y(n932) );
  XOR2xp5r_ASAP7_6t_L U1399 ( .A(n1053), .B(n931), .Y(n1052) );
  OAI22xp5_ASAP7_6t_L U1400 ( .A1(n1054), .A2(n1055), .B1(n1056), .B2(n1057), 
        .Y(n931) );
  NOR2xp5_ASAP7_6t_L U1401 ( .A(n231), .B(n91), .Y(n1053) );
  XOR2xp5r_ASAP7_6t_L U1402 ( .A(n1058), .B(n926), .Y(n927) );
  XOR2xp5r_ASAP7_6t_L U1403 ( .A(n917), .B(n921), .Y(n926) );
  OAI22xp5_ASAP7_6t_L U1404 ( .A1(n1059), .A2(n1060), .B1(n1061), .B2(n1062), 
        .Y(n921) );
  INVx1_ASAP7_6t_L U1405 ( .A(n1059), .Y(n1061) );
  XOR2xp5r_ASAP7_6t_L U1406 ( .A(n1063), .B(n923), .Y(n917) );
  XOR2xp5r_ASAP7_6t_L U1407 ( .A(n1064), .B(n922), .Y(n923) );
  NOR2xp5_ASAP7_6t_L U1408 ( .A(n236), .B(n212), .Y(n922) );
  INVx1_ASAP7_6t_L U1409 ( .A(b[7]), .Y(n212) );
  NAND2xp5R_ASAP7_6t_L U1410 ( .A(a[12]), .B(b[6]), .Y(n1064) );
  XOR2xp5r_ASAP7_6t_L U1411 ( .A(n1065), .B(n919), .Y(n1063) );
  NOR2xp5_ASAP7_6t_L U1412 ( .A(n355), .B(n104), .Y(n919) );
  INVx1_ASAP7_6t_L U1413 ( .A(a[14]), .Y(n104) );
  NAND2xp5R_ASAP7_6t_L U1414 ( .A(b[5]), .B(a[13]), .Y(n1065) );
  AOI21xp25_ASAP7_6t_L U1415 ( .A1(n1066), .A2(n1067), .B(n1068), .Y(n1058) );
  NOR3x1f_ASAP7_6t_L U1416 ( .A(n1066), .B(n102), .C(n355), .Y(n1068) );
  AO22x1_ASAP7_6t_L U1417 ( .A1(n1069), .A2(n1070), .B1(n1071), .B2(n1072), 
        .Y(n930) );
  AOI21xp25_ASAP7_6t_L U1418 ( .A1(n941), .A2(n942), .B(n1073), .Y(n937) );
  NOR3x1f_ASAP7_6t_L U1419 ( .A(n942), .B(n1074), .C(n1075), .Y(n1073) );
  XOR2xp5r_ASAP7_6t_L U1420 ( .A(n1070), .B(n1076), .Y(n942) );
  XOR2xp5r_ASAP7_6t_L U1421 ( .A(n1077), .B(n1069), .Y(n1076) );
  XOR2xp5r_ASAP7_6t_L U1422 ( .A(n1054), .B(n1055), .Y(n1069) );
  INVx1_ASAP7_6t_L U1423 ( .A(n1078), .Y(n1055) );
  XOR2xp5r_ASAP7_6t_L U1424 ( .A(n1056), .B(n1057), .Y(n1078) );
  NAND2xp5R_ASAP7_6t_L U1425 ( .A(a[14]), .B(b[3]), .Y(n1057) );
  NAND2xp5R_ASAP7_6t_L U1426 ( .A(a[15]), .B(b[2]), .Y(n1056) );
  AOI21xp25_ASAP7_6t_L U1427 ( .A1(n1079), .A2(n1080), .B(n1081), .Y(n1054) );
  NOR2xp5_ASAP7_6t_L U1428 ( .A(n1074), .B(n1075), .Y(n1077) );
  INVx1_ASAP7_6t_L U1429 ( .A(n1082), .Y(n1075) );
  INVx1_ASAP7_6t_L U1430 ( .A(n1071), .Y(n1070) );
  XOR2xp5r_ASAP7_6t_L U1431 ( .A(n1083), .B(n1072), .Y(n1071) );
  XOR2xp5r_ASAP7_6t_L U1432 ( .A(n1066), .B(n1067), .Y(n1072) );
  OAI22xp5_ASAP7_6t_L U1433 ( .A1(n1084), .A2(n1085), .B1(n1086), .B2(n1087), 
        .Y(n1067) );
  INVx1_ASAP7_6t_L U1434 ( .A(n1084), .Y(n1086) );
  XOR2xp5r_ASAP7_6t_L U1435 ( .A(n1059), .B(n1088), .Y(n1066) );
  XOR2xp5r_ASAP7_6t_L U1436 ( .A(n1089), .B(n1060), .Y(n1088) );
  NAND2xp5R_ASAP7_6t_L U1437 ( .A(b[5]), .B(a[12]), .Y(n1060) );
  NOR2xp5_ASAP7_6t_L U1438 ( .A(n102), .B(n355), .Y(n1089) );
  XOR2xp5r_ASAP7_6t_L U1439 ( .A(n1090), .B(n1062), .Y(n1059) );
  NAND2xp5R_ASAP7_6t_L U1440 ( .A(b[7]), .B(a[10]), .Y(n1062) );
  NOR2xp5_ASAP7_6t_L U1441 ( .A(n272), .B(n236), .Y(n1090) );
  AOI21xp25_ASAP7_6t_L U1442 ( .A1(n1091), .A2(n1092), .B(n1093), .Y(n1083) );
  NOR3x1f_ASAP7_6t_L U1443 ( .A(n1091), .B(n242), .C(n355), .Y(n1093) );
  OAI22xp5_ASAP7_6t_L U1444 ( .A1(n1094), .A2(n133), .B1(n131), .B2(n1095), 
        .Y(n941) );
  XOR2xp5r_ASAP7_6t_L U1445 ( .A(n1082), .B(n1074), .Y(n133) );
  OA22x1_ASAP7_6t_L U1446 ( .A1(n179), .A2(n182), .B1(n1096), .B2(n1097), .Y(
        n1074) );
  NAND2xp5R_ASAP7_6t_L U1447 ( .A(b[1]), .B(a[14]), .Y(n182) );
  INVx1_ASAP7_6t_L U1448 ( .A(n1096), .Y(n179) );
  XOR2xp5r_ASAP7_6t_L U1449 ( .A(n1097), .B(n1098), .Y(n1096) );
  NAND2xp5R_ASAP7_6t_L U1450 ( .A(b[2]), .B(a[13]), .Y(n1098) );
  NAND2xp5R_ASAP7_6t_L U1451 ( .A(b[3]), .B(a[12]), .Y(n1097) );
  O2A1O1Ixp33_ASAP7_6t_L U1452 ( .A1(n91), .A2(n93), .B(n1080), .C(n1081), .Y(
        n1082) );
  NOR3x1f_ASAP7_6t_L U1453 ( .A(n91), .B(n1080), .C(n93), .Y(n1081) );
  XOR2xp5r_ASAP7_6t_L U1454 ( .A(n1099), .B(n1079), .Y(n1080) );
  NOR2xp5_ASAP7_6t_L U1455 ( .A(n102), .B(n231), .Y(n1079) );
  INVx1_ASAP7_6t_L U1456 ( .A(b[3]), .Y(n231) );
  INVx1_ASAP7_6t_L U1457 ( .A(a[13]), .Y(n102) );
  NAND2xp5R_ASAP7_6t_L U1458 ( .A(b[2]), .B(a[14]), .Y(n1099) );
  INVx1_ASAP7_6t_L U1459 ( .A(b[1]), .Y(n93) );
  INVx1_ASAP7_6t_L U1460 ( .A(a[15]), .Y(n91) );
  INVx1_ASAP7_6t_L U1461 ( .A(n131), .Y(n1094) );
  XOR2xp5r_ASAP7_6t_L U1462 ( .A(n1100), .B(n1095), .Y(n131) );
  INVx1_ASAP7_6t_L U1463 ( .A(n1101), .Y(n1095) );
  XOR2xp5r_ASAP7_6t_L U1464 ( .A(n1091), .B(n1092), .Y(n1101) );
  OAI22xp5_ASAP7_6t_L U1465 ( .A1(n1102), .A2(n1103), .B1(n1104), .B2(n1105), 
        .Y(n1092) );
  XOR2xp5r_ASAP7_6t_L U1466 ( .A(n1084), .B(n1106), .Y(n1091) );
  XOR2xp5r_ASAP7_6t_L U1467 ( .A(n1107), .B(n1085), .Y(n1106) );
  NAND2xp5R_ASAP7_6t_L U1468 ( .A(a[11]), .B(b[5]), .Y(n1085) );
  NOR2xp5_ASAP7_6t_L U1469 ( .A(n242), .B(n355), .Y(n1107) );
  INVx1_ASAP7_6t_L U1470 ( .A(a[12]), .Y(n242) );
  XOR2xp5r_ASAP7_6t_L U1471 ( .A(n1108), .B(n1087), .Y(n1084) );
  NAND2xp5R_ASAP7_6t_L U1472 ( .A(b[7]), .B(a[9]), .Y(n1087) );
  NOR2xp5_ASAP7_6t_L U1473 ( .A(n272), .B(n232), .Y(n1108) );
  AOI21xp25_ASAP7_6t_L U1474 ( .A1(n177), .A2(n178), .B(n1109), .Y(n1100) );
  NOR3x1f_ASAP7_6t_L U1475 ( .A(n177), .B(n355), .C(n236), .Y(n1109) );
  INVx1_ASAP7_6t_L U1476 ( .A(a[11]), .Y(n236) );
  AO21x1_ASAP7_6t_L U1477 ( .A1(n1110), .A2(n233), .B(n1111), .Y(n178) );
  NOR3x1f_ASAP7_6t_L U1478 ( .A(n233), .B(n232), .C(n355), .Y(n1111) );
  INVx1_ASAP7_6t_L U1479 ( .A(b[4]), .Y(n355) );
  INVx1_ASAP7_6t_L U1480 ( .A(a[10]), .Y(n232) );
  XOR2xp5r_ASAP7_6t_L U1481 ( .A(n1112), .B(n1110), .Y(n233) );
  NAND2xp5R_ASAP7_6t_L U1482 ( .A(a[9]), .B(b[5]), .Y(n1112) );
  NOR2xp5_ASAP7_6t_L U1483 ( .A(n272), .B(n301), .Y(n1110) );
  INVx1_ASAP7_6t_L U1484 ( .A(a[8]), .Y(n301) );
  XOR2xp5r_ASAP7_6t_L U1485 ( .A(n1113), .B(n1104), .Y(n177) );
  INVx1_ASAP7_6t_L U1486 ( .A(n1102), .Y(n1104) );
  XOR2xp5r_ASAP7_6t_L U1487 ( .A(n1114), .B(n1105), .Y(n1102) );
  NAND2xp5R_ASAP7_6t_L U1488 ( .A(b[7]), .B(a[8]), .Y(n1105) );
  NOR2xp5_ASAP7_6t_L U1489 ( .A(n356), .B(n272), .Y(n1114) );
  INVx1_ASAP7_6t_L U1490 ( .A(b[6]), .Y(n272) );
  INVx1_ASAP7_6t_L U1491 ( .A(a[9]), .Y(n356) );
  XOR2xp5r_ASAP7_6t_L U1492 ( .A(n1115), .B(n1103), .Y(n1113) );
  NAND2xp5R_ASAP7_6t_L U1493 ( .A(a[10]), .B(b[5]), .Y(n1103) );
  NAND2xp5R_ASAP7_6t_L U1494 ( .A(a[11]), .B(b[4]), .Y(n1115) );
endmodule

