
module DADDA_16x16_52 ( a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [31:0] out;
  wire   n35, n36, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1105, n1107, n1109,
         n1111, n1113, n1115, n1117, n1119, n1121, n1123, n1125, n1127, n1129,
         n1131, n1133, n1135, n1136, n1138, n1140, n1142, n1144, n1146, n1148,
         n1150, n1152, n1154, n1156, n1158, n1159, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216;
  wire   [32:1] p;
  wire   [87:59] s;
  wire   [86:59] c;

  FAxp33_ASAP7_6t_L add_146_U1_1 ( .A(s[59]), .B(p[32]), .CI(n35), .CON(n1162), 
        .SN(n1161) );
  FAxp33_ASAP7_6t_L add_146_U1_2 ( .A(n1158), .B(c[59]), .CI(n1159), .CON(
        n1164), .SN(n1163) );
  FAxp33_ASAP7_6t_L add_146_U1_4 ( .A(s[62]), .B(c[61]), .CI(n36), .CON(n1166), 
        .SN(n1165) );
  FAxp33_ASAP7_6t_L add_146_U1_5 ( .A(s[63]), .B(c[62]), .CI(n1154), .CON(
        n1168), .SN(n1167) );
  FAxp33_ASAP7_6t_L add_146_U1_6 ( .A(s[64]), .B(c[63]), .CI(n1152), .CON(
        n1170), .SN(n1169) );
  FAxp33_ASAP7_6t_L add_146_U1_7 ( .A(s[65]), .B(c[64]), .CI(n1150), .CON(
        n1172), .SN(n1171) );
  FAxp33_ASAP7_6t_L add_146_U1_8 ( .A(s[66]), .B(c[65]), .CI(n1148), .CON(
        n1174), .SN(n1173) );
  FAxp33_ASAP7_6t_L add_146_U1_9 ( .A(s[67]), .B(c[66]), .CI(n1146), .CON(
        n1176), .SN(n1175) );
  FAxp33_ASAP7_6t_L add_146_U1_10 ( .A(s[68]), .B(c[67]), .CI(n1144), .CON(
        n1178), .SN(n1177) );
  FAxp33_ASAP7_6t_L add_146_U1_11 ( .A(s[69]), .B(c[68]), .CI(n1142), .CON(
        n1180), .SN(n1179) );
  FAxp33_ASAP7_6t_L add_146_U1_12 ( .A(s[70]), .B(c[69]), .CI(n1140), .CON(
        n1182), .SN(n1181) );
  FAxp33_ASAP7_6t_L add_146_U1_13 ( .A(s[71]), .B(c[70]), .CI(n1138), .CON(
        n1184), .SN(n1183) );
  FAxp33_ASAP7_6t_L add_146_U1_14 ( .A(s[72]), .B(c[71]), .CI(n1136), .CON(
        n1186), .SN(n1185) );
  FAxp33_ASAP7_6t_L add_146_U1_15 ( .A(s[73]), .B(c[72]), .CI(n1133), .CON(
        n1188), .SN(n1187) );
  FAxp33_ASAP7_6t_L add_146_U1_16 ( .A(s[74]), .B(c[73]), .CI(n1131), .CON(
        n1190), .SN(n1189) );
  FAxp33_ASAP7_6t_L add_146_U1_17 ( .A(s[75]), .B(c[74]), .CI(n1129), .CON(
        n1192), .SN(n1191) );
  FAxp33_ASAP7_6t_L add_146_U1_18 ( .A(s[76]), .B(c[75]), .CI(n1127), .CON(
        n1194), .SN(n1193) );
  FAxp33_ASAP7_6t_L add_146_U1_19 ( .A(s[77]), .B(c[76]), .CI(n1125), .CON(
        n1196), .SN(n1195) );
  FAxp33_ASAP7_6t_L add_146_U1_20 ( .A(s[78]), .B(c[77]), .CI(n1123), .CON(
        n1198), .SN(n1197) );
  FAxp33_ASAP7_6t_L add_146_U1_21 ( .A(s[79]), .B(c[78]), .CI(n1121), .CON(
        n1200), .SN(n1199) );
  FAxp33_ASAP7_6t_L add_146_U1_22 ( .A(s[80]), .B(c[79]), .CI(n1119), .CON(
        n1202), .SN(n1201) );
  FAxp33_ASAP7_6t_L add_146_U1_23 ( .A(s[81]), .B(c[80]), .CI(n1117), .CON(
        n1204), .SN(n1203) );
  FAxp33_ASAP7_6t_L add_146_U1_24 ( .A(s[82]), .B(c[81]), .CI(n1115), .CON(
        n1206), .SN(n1205) );
  FAxp33_ASAP7_6t_L add_146_U1_25 ( .A(s[83]), .B(c[82]), .CI(n1113), .CON(
        n1208), .SN(n1207) );
  FAxp33_ASAP7_6t_L add_146_U1_26 ( .A(s[84]), .B(c[83]), .CI(n1111), .CON(
        n1210), .SN(n1209) );
  FAxp33_ASAP7_6t_L add_146_U1_27 ( .A(s[85]), .B(c[84]), .CI(n1109), .CON(
        n1212), .SN(n1211) );
  FAxp33_ASAP7_6t_L add_146_U1_28 ( .A(s[86]), .B(c[85]), .CI(n1107), .CON(
        n1214), .SN(n1213) );
  FAxp33_ASAP7_6t_L add_146_U1_29 ( .A(s[87]), .B(c[86]), .CI(n1105), .CON(
        n1216), .SN(n1215) );
  AND2x2_ASAP7_6t_L U292 ( .A(p[16]), .B(p[1]), .Y(n35) );
  AND2x2_ASAP7_6t_L U293 ( .A(s[61]), .B(n1156), .Y(n36) );
  XOR2xp5r_ASAP7_6t_L U294 ( .A(p[1]), .B(p[16]), .Y(out[1]) );
  XOR2xp5r_ASAP7_6t_L U295 ( .A(n1156), .B(s[61]), .Y(out[4]) );
  XOR2xp5r_ASAP7_6t_L U296 ( .A(n1135), .B(n1103), .Y(out[31]) );
  XOR2xp5r_ASAP7_6t_L U297 ( .A(n40), .B(n41), .Y(s[87]) );
  XOR2xp5r_ASAP7_6t_L U298 ( .A(n42), .B(n43), .Y(s[86]) );
  XOR2xp5r_ASAP7_6t_L U299 ( .A(n44), .B(n45), .Y(s[85]) );
  XOR2xp5r_ASAP7_6t_L U300 ( .A(n46), .B(n47), .Y(s[84]) );
  XOR2xp5r_ASAP7_6t_L U301 ( .A(n48), .B(n49), .Y(s[83]) );
  XOR2xp5r_ASAP7_6t_L U302 ( .A(n50), .B(n51), .Y(s[82]) );
  XOR2xp5r_ASAP7_6t_L U303 ( .A(n52), .B(n53), .Y(s[81]) );
  XOR2xp5r_ASAP7_6t_L U304 ( .A(n54), .B(n55), .Y(s[80]) );
  XOR2xp5r_ASAP7_6t_L U305 ( .A(n56), .B(n57), .Y(s[79]) );
  XOR2xp5r_ASAP7_6t_L U306 ( .A(n58), .B(n59), .Y(s[78]) );
  XOR2xp5r_ASAP7_6t_L U307 ( .A(n60), .B(n61), .Y(s[77]) );
  XOR2xp5r_ASAP7_6t_L U308 ( .A(n62), .B(n63), .Y(s[76]) );
  XOR2xp5r_ASAP7_6t_L U309 ( .A(n64), .B(n65), .Y(s[75]) );
  XOR2xp5r_ASAP7_6t_L U310 ( .A(n66), .B(n67), .Y(s[74]) );
  XOR2xp5r_ASAP7_6t_L U311 ( .A(n68), .B(n69), .Y(s[73]) );
  XOR2xp5r_ASAP7_6t_L U312 ( .A(n70), .B(n71), .Y(s[72]) );
  XOR2xp5r_ASAP7_6t_L U313 ( .A(n72), .B(n73), .Y(s[71]) );
  XOR2xp5r_ASAP7_6t_L U314 ( .A(n74), .B(n75), .Y(s[70]) );
  XOR2xp5r_ASAP7_6t_L U315 ( .A(n76), .B(n77), .Y(s[69]) );
  XOR2xp5r_ASAP7_6t_L U316 ( .A(n78), .B(n79), .Y(s[68]) );
  XOR2xp5r_ASAP7_6t_L U317 ( .A(n80), .B(n81), .Y(s[67]) );
  XOR2xp5r_ASAP7_6t_L U318 ( .A(n82), .B(n83), .Y(s[66]) );
  XOR2xp5r_ASAP7_6t_L U319 ( .A(n84), .B(n85), .Y(s[65]) );
  XOR2xp5r_ASAP7_6t_L U320 ( .A(n86), .B(n87), .Y(s[64]) );
  XOR2xp5r_ASAP7_6t_L U321 ( .A(n88), .B(n89), .Y(s[63]) );
  XOR2xp5r_ASAP7_6t_L U322 ( .A(n90), .B(n91), .Y(s[62]) );
  XOR2xp5r_ASAP7_6t_L U323 ( .A(n92), .B(n93), .Y(s[61]) );
  XOR2xp5r_ASAP7_6t_L U324 ( .A(n94), .B(n95), .Y(s[59]) );
  NAND2xp5R_ASAP7_6t_L U325 ( .A(b[1]), .B(a[1]), .Y(n94) );
  NOR2xp5_ASAP7_6t_L U326 ( .A(n96), .B(n97), .Y(p[32]) );
  NOR2xp5_ASAP7_6t_L U327 ( .A(n98), .B(n99), .Y(p[1]) );
  NOR2xp5_ASAP7_6t_L U328 ( .A(n100), .B(n97), .Y(p[16]) );
  NOR2xp5_ASAP7_6t_L U329 ( .A(n98), .B(n97), .Y(out[0]) );
  INVx1_ASAP7_6t_L U330 ( .A(n1216), .Y(n1103) );
  INVx1_ASAP7_6t_L U331 ( .A(n1215), .Y(out[30]) );
  INVx1_ASAP7_6t_L U332 ( .A(n1214), .Y(n1105) );
  INVx1_ASAP7_6t_L U333 ( .A(n1213), .Y(out[29]) );
  INVx1_ASAP7_6t_L U334 ( .A(n1212), .Y(n1107) );
  INVx1_ASAP7_6t_L U335 ( .A(n1211), .Y(out[28]) );
  INVx1_ASAP7_6t_L U336 ( .A(n1210), .Y(n1109) );
  INVx1_ASAP7_6t_L U337 ( .A(n1209), .Y(out[27]) );
  INVx1_ASAP7_6t_L U338 ( .A(n1208), .Y(n1111) );
  INVx1_ASAP7_6t_L U339 ( .A(n1207), .Y(out[26]) );
  INVx1_ASAP7_6t_L U340 ( .A(n1206), .Y(n1113) );
  INVx1_ASAP7_6t_L U341 ( .A(n1205), .Y(out[25]) );
  INVx1_ASAP7_6t_L U342 ( .A(n1204), .Y(n1115) );
  INVx1_ASAP7_6t_L U343 ( .A(n1203), .Y(out[24]) );
  INVx1_ASAP7_6t_L U344 ( .A(n1202), .Y(n1117) );
  INVx1_ASAP7_6t_L U345 ( .A(n1201), .Y(out[23]) );
  INVx1_ASAP7_6t_L U346 ( .A(n1200), .Y(n1119) );
  INVx1_ASAP7_6t_L U347 ( .A(n1199), .Y(out[22]) );
  INVx1_ASAP7_6t_L U348 ( .A(n1198), .Y(n1121) );
  INVx1_ASAP7_6t_L U349 ( .A(n1197), .Y(out[21]) );
  INVx1_ASAP7_6t_L U350 ( .A(n1196), .Y(n1123) );
  INVx1_ASAP7_6t_L U351 ( .A(n1195), .Y(out[20]) );
  INVx1_ASAP7_6t_L U352 ( .A(n1194), .Y(n1125) );
  INVx1_ASAP7_6t_L U353 ( .A(n1193), .Y(out[19]) );
  INVx1_ASAP7_6t_L U354 ( .A(n1192), .Y(n1127) );
  INVx1_ASAP7_6t_L U355 ( .A(n1191), .Y(out[18]) );
  INVx1_ASAP7_6t_L U356 ( .A(n1190), .Y(n1129) );
  INVx1_ASAP7_6t_L U357 ( .A(n1189), .Y(out[17]) );
  INVx1_ASAP7_6t_L U358 ( .A(n1188), .Y(n1131) );
  INVx1_ASAP7_6t_L U359 ( .A(n1187), .Y(out[16]) );
  INVx1_ASAP7_6t_L U360 ( .A(n1186), .Y(n1133) );
  INVx1_ASAP7_6t_L U361 ( .A(n1185), .Y(out[15]) );
  OAI22xp5_ASAP7_6t_L U362 ( .A1(n41), .A2(n40), .B1(n101), .B2(n102), .Y(
        n1135) );
  OAI211xp33_ASAP7_6t_L U363 ( .A1(n101), .A2(n102), .B(b[15]), .C(a[15]), .Y(
        n41) );
  INVx1_ASAP7_6t_L U364 ( .A(n1184), .Y(n1136) );
  INVx1_ASAP7_6t_L U365 ( .A(n1183), .Y(out[14]) );
  INVx1_ASAP7_6t_L U366 ( .A(n1182), .Y(n1138) );
  INVx1_ASAP7_6t_L U367 ( .A(n1181), .Y(out[13]) );
  INVx1_ASAP7_6t_L U368 ( .A(n1180), .Y(n1140) );
  INVx1_ASAP7_6t_L U369 ( .A(n1179), .Y(out[12]) );
  INVx1_ASAP7_6t_L U370 ( .A(n1178), .Y(n1142) );
  INVx1_ASAP7_6t_L U371 ( .A(n1177), .Y(out[11]) );
  INVx1_ASAP7_6t_L U372 ( .A(n1176), .Y(n1144) );
  INVx1_ASAP7_6t_L U373 ( .A(n1175), .Y(out[10]) );
  INVx1_ASAP7_6t_L U374 ( .A(n1174), .Y(n1146) );
  INVx1_ASAP7_6t_L U375 ( .A(n1173), .Y(out[9]) );
  INVx1_ASAP7_6t_L U376 ( .A(n1172), .Y(n1148) );
  INVx1_ASAP7_6t_L U377 ( .A(n1171), .Y(out[8]) );
  INVx1_ASAP7_6t_L U378 ( .A(n1170), .Y(n1150) );
  INVx1_ASAP7_6t_L U379 ( .A(n1169), .Y(out[7]) );
  INVx1_ASAP7_6t_L U380 ( .A(n1168), .Y(n1152) );
  INVx1_ASAP7_6t_L U381 ( .A(n1167), .Y(out[6]) );
  INVx1_ASAP7_6t_L U382 ( .A(n1166), .Y(n1154) );
  INVx1_ASAP7_6t_L U383 ( .A(n1165), .Y(out[5]) );
  INVx1_ASAP7_6t_L U384 ( .A(n1164), .Y(n1156) );
  INVx1_ASAP7_6t_L U385 ( .A(n1163), .Y(out[3]) );
  INVx1_ASAP7_6t_L U386 ( .A(n1162), .Y(n1159) );
  INVx1_ASAP7_6t_L U387 ( .A(n1161), .Y(out[2]) );
  NOR2xp5_ASAP7_6t_L U388 ( .A(n43), .B(n42), .Y(c[86]) );
  OAI21xp25_ASAP7_6t_L U389 ( .A1(n102), .A2(n103), .B(n40), .Y(n42) );
  NAND2xp5R_ASAP7_6t_L U390 ( .A(n102), .B(n103), .Y(n40) );
  OAI21xp25_ASAP7_6t_L U391 ( .A1(n104), .A2(n105), .B(n106), .Y(n103) );
  XOR2xp5r_ASAP7_6t_L U392 ( .A(n107), .B(n101), .Y(n102) );
  NAND2xp5R_ASAP7_6t_L U393 ( .A(a[14]), .B(b[15]), .Y(n101) );
  NAND2xp5R_ASAP7_6t_L U394 ( .A(b[14]), .B(a[15]), .Y(n107) );
  NOR2xp5_ASAP7_6t_L U395 ( .A(n45), .B(n44), .Y(c[85]) );
  OAI21xp25_ASAP7_6t_L U396 ( .A1(n108), .A2(n109), .B(n43), .Y(n44) );
  NAND2xp5R_ASAP7_6t_L U397 ( .A(n108), .B(n109), .Y(n43) );
  OR2x2_ASAP7_6t_L U398 ( .A(n110), .B(n111), .Y(n109) );
  NOR3x1f_ASAP7_6t_L U399 ( .A(n112), .B(n113), .C(n114), .Y(n111) );
  NOR3x1f_ASAP7_6t_L U400 ( .A(n115), .B(n116), .C(n117), .Y(n110) );
  INVx1_ASAP7_6t_L U401 ( .A(n112), .Y(n115) );
  INVx1_ASAP7_6t_L U402 ( .A(n118), .Y(n108) );
  A2O1A1Ixp33_ASAP7_6t_L U403 ( .A1(b[13]), .A2(a[15]), .B(n105), .C(n106), 
        .Y(n118) );
  NAND3xp33R_ASAP7_6t_L U404 ( .A(b[13]), .B(n105), .C(a[15]), .Y(n106) );
  XOR2xp5r_ASAP7_6t_L U405 ( .A(n104), .B(n119), .Y(n105) );
  NAND2xp5R_ASAP7_6t_L U406 ( .A(b[14]), .B(a[14]), .Y(n119) );
  NAND2xp5R_ASAP7_6t_L U407 ( .A(b[15]), .B(a[13]), .Y(n104) );
  OA22x1_ASAP7_6t_L U408 ( .A1(n120), .A2(n121), .B1(n122), .B2(n123), .Y(n45)
         );
  AO21x1_ASAP7_6t_L U409 ( .A1(n46), .A2(n47), .B(n124), .Y(c[84]) );
  NOR3x1f_ASAP7_6t_L U410 ( .A(n47), .B(n125), .C(n126), .Y(n124) );
  XOR2xp5r_ASAP7_6t_L U411 ( .A(n127), .B(n123), .Y(n47) );
  AOI21xp25_ASAP7_6t_L U412 ( .A1(n128), .A2(n129), .B(n130), .Y(n123) );
  NOR3x1f_ASAP7_6t_L U413 ( .A(n129), .B(n131), .C(n126), .Y(n130) );
  XOR2xp5r_ASAP7_6t_L U414 ( .A(n132), .B(n122), .Y(n127) );
  INVx1_ASAP7_6t_L U415 ( .A(n120), .Y(n122) );
  XOR2xp5r_ASAP7_6t_L U416 ( .A(n133), .B(n112), .Y(n120) );
  XOR2xp5r_ASAP7_6t_L U417 ( .A(n134), .B(n135), .Y(n112) );
  NAND2xp5R_ASAP7_6t_L U418 ( .A(a[12]), .B(b[15]), .Y(n135) );
  AOI22xp25_ASAP7_6t_L U419 ( .A1(n136), .A2(n137), .B1(n138), .B2(n139), .Y(
        n134) );
  XOR2xp5r_ASAP7_6t_L U420 ( .A(n140), .B(n121), .Y(n133) );
  NAND2xp5R_ASAP7_6t_L U421 ( .A(b[13]), .B(a[14]), .Y(n121) );
  NAND2xp5R_ASAP7_6t_L U422 ( .A(b[14]), .B(a[13]), .Y(n140) );
  NOR2xp5_ASAP7_6t_L U423 ( .A(n125), .B(n126), .Y(n132) );
  OAI22xp5_ASAP7_6t_L U424 ( .A1(n141), .A2(n142), .B1(n143), .B2(n144), .Y(
        n46) );
  AO21x1_ASAP7_6t_L U425 ( .A1(n48), .A2(n49), .B(n145), .Y(c[83]) );
  NOR3x1f_ASAP7_6t_L U426 ( .A(n48), .B(n125), .C(n146), .Y(n145) );
  AO21x1_ASAP7_6t_L U427 ( .A1(n147), .A2(n148), .B(n149), .Y(n49) );
  NOR3x1f_ASAP7_6t_L U428 ( .A(n147), .B(n131), .C(n146), .Y(n149) );
  XOR2xp5r_ASAP7_6t_L U429 ( .A(n141), .B(n150), .Y(n48) );
  XOR2xp5r_ASAP7_6t_L U430 ( .A(n151), .B(n142), .Y(n150) );
  INVx1_ASAP7_6t_L U431 ( .A(n144), .Y(n142) );
  XOR2xp5r_ASAP7_6t_L U432 ( .A(n129), .B(n152), .Y(n144) );
  XOR2xp5r_ASAP7_6t_L U433 ( .A(n153), .B(n143), .Y(n152) );
  AOI22xp25_ASAP7_6t_L U434 ( .A1(n154), .A2(n155), .B1(n156), .B2(n157), .Y(
        n143) );
  NOR2xp5_ASAP7_6t_L U435 ( .A(n131), .B(n126), .Y(n153) );
  XOR2xp5r_ASAP7_6t_L U436 ( .A(n158), .B(n128), .Y(n129) );
  XOR2xp5r_ASAP7_6t_L U437 ( .A(n139), .B(n138), .Y(n128) );
  NOR2xp5_ASAP7_6t_L U438 ( .A(n159), .B(n116), .Y(n138) );
  XOR2xp5r_ASAP7_6t_L U439 ( .A(n137), .B(n136), .Y(n139) );
  NOR2xp5_ASAP7_6t_L U440 ( .A(n114), .B(n117), .Y(n136) );
  NOR2xp5_ASAP7_6t_L U441 ( .A(n160), .B(n113), .Y(n137) );
  AOI22xp25_ASAP7_6t_L U442 ( .A1(n161), .A2(n162), .B1(n163), .B2(n164), .Y(
        n158) );
  NOR2xp5_ASAP7_6t_L U443 ( .A(n125), .B(n146), .Y(n151) );
  AOI22xp25_ASAP7_6t_L U444 ( .A1(n165), .A2(n166), .B1(n167), .B2(n168), .Y(
        n141) );
  AO21x1_ASAP7_6t_L U445 ( .A1(n50), .A2(n51), .B(n169), .Y(c[82]) );
  NOR3x1f_ASAP7_6t_L U446 ( .A(n50), .B(n125), .C(n170), .Y(n169) );
  OAI22xp5_ASAP7_6t_L U447 ( .A1(n171), .A2(n172), .B1(n173), .B2(n174), .Y(
        n51) );
  XOR2xp5r_ASAP7_6t_L U448 ( .A(n175), .B(n148), .Y(n50) );
  AO21x1_ASAP7_6t_L U449 ( .A1(n176), .A2(n177), .B(n178), .Y(n148) );
  NOR3x1f_ASAP7_6t_L U450 ( .A(n177), .B(n131), .C(n170), .Y(n178) );
  XOR2xp5r_ASAP7_6t_L U451 ( .A(n179), .B(n147), .Y(n175) );
  XOR2xp5r_ASAP7_6t_L U452 ( .A(n180), .B(n165), .Y(n147) );
  INVx1_ASAP7_6t_L U453 ( .A(n167), .Y(n165) );
  XOR2xp5r_ASAP7_6t_L U454 ( .A(n181), .B(n168), .Y(n167) );
  XOR2xp5r_ASAP7_6t_L U455 ( .A(n164), .B(n163), .Y(n168) );
  AO21x1_ASAP7_6t_L U456 ( .A1(n182), .A2(n183), .B(n184), .Y(n163) );
  NOR3x1f_ASAP7_6t_L U457 ( .A(n183), .B(n159), .C(n160), .Y(n184) );
  XOR2xp5r_ASAP7_6t_L U458 ( .A(n161), .B(n162), .Y(n164) );
  NOR2xp5_ASAP7_6t_L U459 ( .A(n185), .B(n113), .Y(n162) );
  NOR2xp5_ASAP7_6t_L U460 ( .A(n160), .B(n117), .Y(n161) );
  AOI21xp25_ASAP7_6t_L U461 ( .A1(n186), .A2(n187), .B(n188), .Y(n181) );
  NOR3x1f_ASAP7_6t_L U462 ( .A(n186), .B(n116), .C(n146), .Y(n188) );
  XOR2xp5r_ASAP7_6t_L U463 ( .A(n189), .B(n166), .Y(n180) );
  XOR2xp5r_ASAP7_6t_L U464 ( .A(n154), .B(n155), .Y(n166) );
  OAI22xp5_ASAP7_6t_L U465 ( .A1(n190), .A2(n191), .B1(n192), .B2(n193), .Y(
        n155) );
  XOR2xp5r_ASAP7_6t_L U466 ( .A(n157), .B(n156), .Y(n154) );
  NOR2xp5_ASAP7_6t_L U467 ( .A(n114), .B(n159), .Y(n156) );
  NOR2xp5_ASAP7_6t_L U468 ( .A(n126), .B(n116), .Y(n157) );
  NOR2xp5_ASAP7_6t_L U469 ( .A(n131), .B(n146), .Y(n189) );
  NOR2xp5_ASAP7_6t_L U470 ( .A(n125), .B(n170), .Y(n179) );
  AO21x1_ASAP7_6t_L U471 ( .A1(n53), .A2(n52), .B(n194), .Y(c[81]) );
  NOR3x1f_ASAP7_6t_L U472 ( .A(n52), .B(n125), .C(n195), .Y(n194) );
  XOR2xp5r_ASAP7_6t_L U473 ( .A(n196), .B(n174), .Y(n52) );
  AOI22xp25_ASAP7_6t_L U474 ( .A1(n197), .A2(n198), .B1(n199), .B2(n200), .Y(
        n174) );
  XOR2xp5r_ASAP7_6t_L U475 ( .A(n201), .B(n173), .Y(n196) );
  INVx1_ASAP7_6t_L U476 ( .A(n172), .Y(n173) );
  XOR2xp5r_ASAP7_6t_L U477 ( .A(n202), .B(n177), .Y(n172) );
  XOR2xp5r_ASAP7_6t_L U478 ( .A(n203), .B(n176), .Y(n177) );
  XOR2xp5r_ASAP7_6t_L U479 ( .A(n187), .B(n186), .Y(n176) );
  XOR2xp5r_ASAP7_6t_L U480 ( .A(n204), .B(n190), .Y(n186) );
  AOI21xp25_ASAP7_6t_L U481 ( .A1(n205), .A2(n206), .B(n207), .Y(n190) );
  NOR3x1f_ASAP7_6t_L U482 ( .A(n206), .B(n159), .C(n185), .Y(n207) );
  XOR2xp5r_ASAP7_6t_L U483 ( .A(n208), .B(n191), .Y(n204) );
  INVx1_ASAP7_6t_L U484 ( .A(n192), .Y(n191) );
  XOR2xp5r_ASAP7_6t_L U485 ( .A(n183), .B(n209), .Y(n192) );
  XOR2xp5r_ASAP7_6t_L U486 ( .A(n210), .B(n193), .Y(n209) );
  NAND2xp5R_ASAP7_6t_L U487 ( .A(b[12]), .B(a[12]), .Y(n193) );
  NOR2xp5_ASAP7_6t_L U488 ( .A(n159), .B(n160), .Y(n210) );
  XOR2xp5r_ASAP7_6t_L U489 ( .A(n211), .B(n182), .Y(n183) );
  NOR2xp5_ASAP7_6t_L U490 ( .A(n212), .B(n113), .Y(n182) );
  NAND2xp5R_ASAP7_6t_L U491 ( .A(b[14]), .B(a[10]), .Y(n211) );
  NOR2xp5_ASAP7_6t_L U492 ( .A(n116), .B(n146), .Y(n208) );
  OAI22xp5_ASAP7_6t_L U493 ( .A1(n213), .A2(n214), .B1(n215), .B2(n216), .Y(
        n187) );
  AOI21xp25_ASAP7_6t_L U494 ( .A1(n217), .A2(n218), .B(n219), .Y(n203) );
  NOR3x1f_ASAP7_6t_L U495 ( .A(n217), .B(n114), .C(n146), .Y(n219) );
  XOR2xp5r_ASAP7_6t_L U496 ( .A(n171), .B(n220), .Y(n202) );
  NOR2xp5_ASAP7_6t_L U497 ( .A(n131), .B(n170), .Y(n220) );
  AOI22xp25_ASAP7_6t_L U498 ( .A1(n221), .A2(n222), .B1(n223), .B2(n224), .Y(
        n171) );
  NOR2xp5_ASAP7_6t_L U499 ( .A(n125), .B(n195), .Y(n201) );
  OAI22xp5_ASAP7_6t_L U500 ( .A1(n225), .A2(n226), .B1(n227), .B2(n228), .Y(
        n53) );
  OAI22xp5_ASAP7_6t_L U501 ( .A1(n54), .A2(n55), .B1(n229), .B2(n230), .Y(
        c[80]) );
  INVx1_ASAP7_6t_L U502 ( .A(n230), .Y(n55) );
  XOR2xp5r_ASAP7_6t_L U503 ( .A(n231), .B(n228), .Y(n230) );
  AOI22xp25_ASAP7_6t_L U504 ( .A1(n232), .A2(n233), .B1(n234), .B2(n235), .Y(
        n228) );
  INVx1_ASAP7_6t_L U505 ( .A(n234), .Y(n232) );
  XOR2xp5r_ASAP7_6t_L U506 ( .A(n229), .B(n226), .Y(n231) );
  INVx1_ASAP7_6t_L U507 ( .A(n227), .Y(n226) );
  XOR2xp5r_ASAP7_6t_L U508 ( .A(n198), .B(n236), .Y(n227) );
  XOR2xp5r_ASAP7_6t_L U509 ( .A(n225), .B(n197), .Y(n236) );
  INVx1_ASAP7_6t_L U510 ( .A(n199), .Y(n197) );
  XOR2xp5r_ASAP7_6t_L U511 ( .A(n237), .B(n200), .Y(n199) );
  XOR2xp5r_ASAP7_6t_L U512 ( .A(n217), .B(n218), .Y(n200) );
  OAI22xp5_ASAP7_6t_L U513 ( .A1(n238), .A2(n239), .B1(n240), .B2(n241), .Y(
        n218) );
  XOR2xp5r_ASAP7_6t_L U514 ( .A(n242), .B(n213), .Y(n217) );
  AOI21xp25_ASAP7_6t_L U515 ( .A1(n243), .A2(n244), .B(n245), .Y(n213) );
  NOR3x1f_ASAP7_6t_L U516 ( .A(n244), .B(n159), .C(n212), .Y(n245) );
  XOR2xp5r_ASAP7_6t_L U517 ( .A(n246), .B(n214), .Y(n242) );
  INVx1_ASAP7_6t_L U518 ( .A(n215), .Y(n214) );
  XOR2xp5r_ASAP7_6t_L U519 ( .A(n206), .B(n247), .Y(n215) );
  XOR2xp5r_ASAP7_6t_L U520 ( .A(n248), .B(n216), .Y(n247) );
  NAND2xp5R_ASAP7_6t_L U521 ( .A(b[12]), .B(a[11]), .Y(n216) );
  NOR2xp5_ASAP7_6t_L U522 ( .A(n159), .B(n185), .Y(n248) );
  XOR2xp5r_ASAP7_6t_L U523 ( .A(n205), .B(n249), .Y(n206) );
  NAND2xp5R_ASAP7_6t_L U524 ( .A(a[9]), .B(b[14]), .Y(n249) );
  NOR2xp5_ASAP7_6t_L U525 ( .A(n250), .B(n113), .Y(n205) );
  NOR2xp5_ASAP7_6t_L U526 ( .A(n114), .B(n146), .Y(n246) );
  AOI21xp25_ASAP7_6t_L U527 ( .A1(n251), .A2(n252), .B(n253), .Y(n237) );
  NOR3x1f_ASAP7_6t_L U528 ( .A(n251), .B(n160), .C(n146), .Y(n253) );
  AOI22xp25_ASAP7_6t_L U529 ( .A1(n254), .A2(n255), .B1(n256), .B2(n257), .Y(
        n225) );
  XOR2xp5r_ASAP7_6t_L U530 ( .A(n221), .B(n222), .Y(n198) );
  NOR2xp5_ASAP7_6t_L U531 ( .A(n258), .B(n125), .Y(n222) );
  XOR2xp5r_ASAP7_6t_L U532 ( .A(n223), .B(n224), .Y(n221) );
  NOR2xp5_ASAP7_6t_L U533 ( .A(n195), .B(n131), .Y(n224) );
  NOR2xp5_ASAP7_6t_L U534 ( .A(n170), .B(n116), .Y(n223) );
  AOI22xp25_ASAP7_6t_L U535 ( .A1(n259), .A2(n260), .B1(n261), .B2(n262), .Y(
        n229) );
  OA22x1_ASAP7_6t_L U536 ( .A1(n263), .A2(n264), .B1(n265), .B2(n266), .Y(n54)
         );
  INVx1_ASAP7_6t_L U537 ( .A(n265), .Y(n264) );
  OAI22xp5_ASAP7_6t_L U538 ( .A1(n57), .A2(n56), .B1(n267), .B2(n268), .Y(
        c[79]) );
  INVx1_ASAP7_6t_L U539 ( .A(n267), .Y(n56) );
  XOR2xp5r_ASAP7_6t_L U540 ( .A(n263), .B(n269), .Y(n267) );
  XOR2xp5r_ASAP7_6t_L U541 ( .A(n268), .B(n265), .Y(n269) );
  XOR2xp5r_ASAP7_6t_L U542 ( .A(n266), .B(n270), .Y(n265) );
  XOR2xp5r_ASAP7_6t_L U543 ( .A(n233), .B(n234), .Y(n270) );
  XOR2xp5r_ASAP7_6t_L U544 ( .A(n271), .B(n235), .Y(n234) );
  XOR2xp5r_ASAP7_6t_L U545 ( .A(n251), .B(n252), .Y(n235) );
  OAI22xp5_ASAP7_6t_L U546 ( .A1(n272), .A2(n273), .B1(n274), .B2(n275), .Y(
        n252) );
  XOR2xp5r_ASAP7_6t_L U547 ( .A(n238), .B(n276), .Y(n251) );
  XOR2xp5r_ASAP7_6t_L U548 ( .A(n240), .B(n277), .Y(n276) );
  NAND2xp5R_ASAP7_6t_L U549 ( .A(b[11]), .B(a[11]), .Y(n277) );
  INVx1_ASAP7_6t_L U550 ( .A(n239), .Y(n240) );
  XOR2xp5r_ASAP7_6t_L U551 ( .A(n278), .B(n244), .Y(n239) );
  XOR2xp5r_ASAP7_6t_L U552 ( .A(n279), .B(n243), .Y(n244) );
  NOR2xp5_ASAP7_6t_L U553 ( .A(n280), .B(n113), .Y(n243) );
  NAND2xp5R_ASAP7_6t_L U554 ( .A(b[14]), .B(a[8]), .Y(n279) );
  XOR2xp5r_ASAP7_6t_L U555 ( .A(n281), .B(n241), .Y(n278) );
  NAND2xp5R_ASAP7_6t_L U556 ( .A(b[12]), .B(a[10]), .Y(n241) );
  NAND2xp5R_ASAP7_6t_L U557 ( .A(a[9]), .B(b[13]), .Y(n281) );
  NOR2xp5_ASAP7_6t_L U558 ( .A(n282), .B(n283), .Y(n238) );
  NOR3x1f_ASAP7_6t_L U559 ( .A(n284), .B(n113), .C(n285), .Y(n283) );
  NOR3x1f_ASAP7_6t_L U560 ( .A(n286), .B(n117), .C(n280), .Y(n282) );
  INVx1_ASAP7_6t_L U561 ( .A(n284), .Y(n286) );
  AOI21xp25_ASAP7_6t_L U562 ( .A1(n287), .A2(n288), .B(n289), .Y(n271) );
  NOR3x1f_ASAP7_6t_L U563 ( .A(n288), .B(n212), .C(n126), .Y(n289) );
  XOR2xp5r_ASAP7_6t_L U564 ( .A(n254), .B(n255), .Y(n233) );
  AO21x1_ASAP7_6t_L U565 ( .A1(n290), .A2(n291), .B(n292), .Y(n255) );
  NOR3x1f_ASAP7_6t_L U566 ( .A(n291), .B(n114), .C(n195), .Y(n292) );
  XOR2xp5r_ASAP7_6t_L U567 ( .A(n257), .B(n256), .Y(n254) );
  NOR2xp5_ASAP7_6t_L U568 ( .A(n170), .B(n114), .Y(n256) );
  NOR2xp5_ASAP7_6t_L U569 ( .A(n195), .B(n116), .Y(n257) );
  AOI21xp25_ASAP7_6t_L U570 ( .A1(n293), .A2(n294), .B(n295), .Y(n266) );
  NOR3x1f_ASAP7_6t_L U571 ( .A(n293), .B(n131), .C(n296), .Y(n295) );
  XOR2xp5r_ASAP7_6t_L U572 ( .A(n297), .B(n260), .Y(n268) );
  OAI22xp5_ASAP7_6t_L U573 ( .A1(n298), .A2(n299), .B1(n300), .B2(n301), .Y(
        n260) );
  INVx1_ASAP7_6t_L U574 ( .A(n299), .Y(n300) );
  INVx1_ASAP7_6t_L U575 ( .A(n259), .Y(n297) );
  XOR2xp5r_ASAP7_6t_L U576 ( .A(n261), .B(n262), .Y(n259) );
  NOR2xp5_ASAP7_6t_L U577 ( .A(n296), .B(n125), .Y(n262) );
  NOR2xp5_ASAP7_6t_L U578 ( .A(n258), .B(n131), .Y(n261) );
  AOI22xp25_ASAP7_6t_L U579 ( .A1(n302), .A2(n303), .B1(n304), .B2(n305), .Y(
        n263) );
  INVx1_ASAP7_6t_L U580 ( .A(n303), .Y(n304) );
  AOI22xp25_ASAP7_6t_L U581 ( .A1(n306), .A2(n307), .B1(n308), .B2(n309), .Y(
        n57) );
  AO21x1_ASAP7_6t_L U582 ( .A1(n59), .A2(n58), .B(n310), .Y(c[78]) );
  NOR3x1f_ASAP7_6t_L U583 ( .A(n58), .B(n125), .C(n311), .Y(n310) );
  XOR2xp5r_ASAP7_6t_L U584 ( .A(n309), .B(n312), .Y(n58) );
  XOR2xp5r_ASAP7_6t_L U585 ( .A(n313), .B(n308), .Y(n312) );
  INVx1_ASAP7_6t_L U586 ( .A(n307), .Y(n308) );
  XOR2xp5r_ASAP7_6t_L U587 ( .A(n306), .B(n314), .Y(n307) );
  XOR2xp5r_ASAP7_6t_L U588 ( .A(n305), .B(n303), .Y(n314) );
  XOR2xp5r_ASAP7_6t_L U589 ( .A(n315), .B(n302), .Y(n303) );
  XOR2xp5r_ASAP7_6t_L U590 ( .A(n287), .B(n288), .Y(n302) );
  XOR2xp5r_ASAP7_6t_L U591 ( .A(n316), .B(n275), .Y(n288) );
  AOI21xp25_ASAP7_6t_L U592 ( .A1(n317), .A2(n318), .B(n319), .Y(n275) );
  NOR3x1f_ASAP7_6t_L U593 ( .A(n318), .B(n126), .C(n250), .Y(n319) );
  XOR2xp5r_ASAP7_6t_L U594 ( .A(n320), .B(n274), .Y(n316) );
  INVx1_ASAP7_6t_L U595 ( .A(n272), .Y(n274) );
  XOR2xp5r_ASAP7_6t_L U596 ( .A(n321), .B(n284), .Y(n272) );
  XOR2xp5r_ASAP7_6t_L U597 ( .A(n322), .B(n323), .Y(n284) );
  NAND2xp5R_ASAP7_6t_L U598 ( .A(a[6]), .B(b[15]), .Y(n323) );
  AOI22xp25_ASAP7_6t_L U599 ( .A1(n324), .A2(n325), .B1(n326), .B2(n327), .Y(
        n322) );
  XOR2xp5r_ASAP7_6t_L U600 ( .A(n328), .B(n273), .Y(n321) );
  NAND2xp5R_ASAP7_6t_L U601 ( .A(a[8]), .B(b[13]), .Y(n273) );
  NAND2xp5R_ASAP7_6t_L U602 ( .A(a[7]), .B(b[14]), .Y(n328) );
  NOR2xp5_ASAP7_6t_L U603 ( .A(n212), .B(n126), .Y(n320) );
  OAI22xp5_ASAP7_6t_L U604 ( .A1(n329), .A2(n330), .B1(n331), .B2(n332), .Y(
        n287) );
  INVx1_ASAP7_6t_L U605 ( .A(n333), .Y(n331) );
  AOI21xp25_ASAP7_6t_L U606 ( .A1(n334), .A2(n335), .B(n336), .Y(n315) );
  NOR3x1f_ASAP7_6t_L U607 ( .A(n334), .B(n212), .C(n146), .Y(n336) );
  XOR2xp5r_ASAP7_6t_L U608 ( .A(n293), .B(n294), .Y(n305) );
  OAI22xp5_ASAP7_6t_L U609 ( .A1(n337), .A2(n338), .B1(n339), .B2(n340), .Y(
        n294) );
  INVx1_ASAP7_6t_L U610 ( .A(n338), .Y(n339) );
  XOR2xp5r_ASAP7_6t_L U611 ( .A(n341), .B(n298), .Y(n293) );
  AOI21xp25_ASAP7_6t_L U612 ( .A1(n342), .A2(n343), .B(n344), .Y(n298) );
  NOR3x1f_ASAP7_6t_L U613 ( .A(n343), .B(n114), .C(n258), .Y(n344) );
  XOR2xp5r_ASAP7_6t_L U614 ( .A(n345), .B(n299), .Y(n341) );
  XOR2xp5r_ASAP7_6t_L U615 ( .A(n346), .B(n291), .Y(n299) );
  XOR2xp5r_ASAP7_6t_L U616 ( .A(n347), .B(n290), .Y(n291) );
  NOR2xp5_ASAP7_6t_L U617 ( .A(n146), .B(n185), .Y(n290) );
  NAND2xp5R_ASAP7_6t_L U618 ( .A(a[11]), .B(b[10]), .Y(n347) );
  XOR2xp5r_ASAP7_6t_L U619 ( .A(n348), .B(n301), .Y(n346) );
  NAND2xp5R_ASAP7_6t_L U620 ( .A(b[8]), .B(a[13]), .Y(n301) );
  NAND2xp5R_ASAP7_6t_L U621 ( .A(b[9]), .B(a[12]), .Y(n348) );
  NOR2xp5_ASAP7_6t_L U622 ( .A(n131), .B(n296), .Y(n345) );
  AO21x1_ASAP7_6t_L U623 ( .A1(n349), .A2(n350), .B(n351), .Y(n306) );
  NOR3x1f_ASAP7_6t_L U624 ( .A(n349), .B(n131), .C(n311), .Y(n351) );
  NOR2xp5_ASAP7_6t_L U625 ( .A(n125), .B(n311), .Y(n313) );
  AO22x1_ASAP7_6t_L U626 ( .A1(n352), .A2(n353), .B1(n354), .B2(n355), .Y(n309) );
  OAI22xp5_ASAP7_6t_L U627 ( .A1(n356), .A2(n357), .B1(n358), .B2(n359), .Y(
        n59) );
  INVx1_ASAP7_6t_L U628 ( .A(n357), .Y(n358) );
  AO21x1_ASAP7_6t_L U629 ( .A1(n61), .A2(n60), .B(n360), .Y(c[77]) );
  NOR3x1f_ASAP7_6t_L U630 ( .A(n61), .B(n125), .C(n361), .Y(n360) );
  OAI22xp5_ASAP7_6t_L U631 ( .A1(n362), .A2(n363), .B1(n364), .B2(n365), .Y(
        n60) );
  INVx1_ASAP7_6t_L U632 ( .A(n364), .Y(n363) );
  XOR2xp5r_ASAP7_6t_L U633 ( .A(n356), .B(n366), .Y(n61) );
  XOR2xp5r_ASAP7_6t_L U634 ( .A(n367), .B(n357), .Y(n366) );
  XOR2xp5r_ASAP7_6t_L U635 ( .A(n359), .B(n368), .Y(n357) );
  XOR2xp5r_ASAP7_6t_L U636 ( .A(n353), .B(n352), .Y(n368) );
  INVx1_ASAP7_6t_L U637 ( .A(n354), .Y(n352) );
  AOI22xp25_ASAP7_6t_L U638 ( .A1(n369), .A2(n370), .B1(n371), .B2(n372), .Y(
        n354) );
  XOR2xp5r_ASAP7_6t_L U639 ( .A(n373), .B(n355), .Y(n372) );
  INVx1_ASAP7_6t_L U640 ( .A(n369), .Y(n371) );
  XOR2xp5r_ASAP7_6t_L U641 ( .A(n374), .B(n355), .Y(n370) );
  XOR2xp5r_ASAP7_6t_L U642 ( .A(n334), .B(n335), .Y(n355) );
  OAI22xp5_ASAP7_6t_L U643 ( .A1(n375), .A2(n376), .B1(n377), .B2(n378), .Y(
        n335) );
  INVx1_ASAP7_6t_L U644 ( .A(n376), .Y(n377) );
  XOR2xp5r_ASAP7_6t_L U645 ( .A(n379), .B(n329), .Y(n334) );
  AOI22xp25_ASAP7_6t_L U646 ( .A1(n380), .A2(n381), .B1(n382), .B2(n383), .Y(
        n329) );
  XOR2xp5r_ASAP7_6t_L U647 ( .A(n384), .B(n330), .Y(n379) );
  INVx1_ASAP7_6t_L U648 ( .A(n332), .Y(n330) );
  XOR2xp5r_ASAP7_6t_L U649 ( .A(n318), .B(n385), .Y(n332) );
  XOR2xp5r_ASAP7_6t_L U650 ( .A(n333), .B(n386), .Y(n385) );
  NAND2xp5R_ASAP7_6t_L U651 ( .A(a[8]), .B(b[12]), .Y(n386) );
  OAI22xp5_ASAP7_6t_L U652 ( .A1(n387), .A2(n388), .B1(n389), .B2(n390), .Y(
        n333) );
  XOR2xp5r_ASAP7_6t_L U653 ( .A(n391), .B(n317), .Y(n318) );
  XOR2xp5r_ASAP7_6t_L U654 ( .A(n327), .B(n326), .Y(n317) );
  NOR2xp5_ASAP7_6t_L U655 ( .A(n280), .B(n159), .Y(n326) );
  XOR2xp5r_ASAP7_6t_L U656 ( .A(n324), .B(n325), .Y(n327) );
  NOR2xp5_ASAP7_6t_L U657 ( .A(n392), .B(n113), .Y(n325) );
  NOR2xp5_ASAP7_6t_L U658 ( .A(n285), .B(n117), .Y(n324) );
  AOI22xp25_ASAP7_6t_L U659 ( .A1(n393), .A2(n394), .B1(n395), .B2(n396), .Y(
        n391) );
  NOR2xp5_ASAP7_6t_L U660 ( .A(n212), .B(n146), .Y(n384) );
  XOR2xp5r_ASAP7_6t_L U661 ( .A(n349), .B(n350), .Y(n353) );
  OAI22xp5_ASAP7_6t_L U662 ( .A1(n397), .A2(n398), .B1(n399), .B2(n400), .Y(
        n350) );
  INVx1_ASAP7_6t_L U663 ( .A(n398), .Y(n399) );
  XOR2xp5r_ASAP7_6t_L U664 ( .A(n401), .B(n337), .Y(n349) );
  AOI21xp25_ASAP7_6t_L U665 ( .A1(n402), .A2(n403), .B(n404), .Y(n337) );
  NOR3x1f_ASAP7_6t_L U666 ( .A(n403), .B(n114), .C(n296), .Y(n404) );
  XOR2xp5r_ASAP7_6t_L U667 ( .A(n405), .B(n338), .Y(n401) );
  XOR2xp5r_ASAP7_6t_L U668 ( .A(n406), .B(n343), .Y(n338) );
  XOR2xp5r_ASAP7_6t_L U669 ( .A(n407), .B(n342), .Y(n343) );
  NOR2xp5_ASAP7_6t_L U670 ( .A(n170), .B(n185), .Y(n342) );
  NAND2xp5R_ASAP7_6t_L U671 ( .A(a[11]), .B(b[9]), .Y(n407) );
  XOR2xp5r_ASAP7_6t_L U672 ( .A(n408), .B(n340), .Y(n406) );
  NAND2xp5R_ASAP7_6t_L U673 ( .A(b[7]), .B(a[13]), .Y(n340) );
  NAND2xp5R_ASAP7_6t_L U674 ( .A(b[8]), .B(a[12]), .Y(n408) );
  NOR2xp5_ASAP7_6t_L U675 ( .A(n131), .B(n311), .Y(n405) );
  AOI21xp25_ASAP7_6t_L U676 ( .A1(n409), .A2(n410), .B(n411), .Y(n359) );
  NOR3x1f_ASAP7_6t_L U677 ( .A(n409), .B(n131), .C(n361), .Y(n411) );
  NOR2xp5_ASAP7_6t_L U678 ( .A(n125), .B(n361), .Y(n367) );
  AOI22xp25_ASAP7_6t_L U679 ( .A1(n412), .A2(n413), .B1(n414), .B2(n415), .Y(
        n356) );
  INVx1_ASAP7_6t_L U680 ( .A(n414), .Y(n412) );
  AO21x1_ASAP7_6t_L U681 ( .A1(n62), .A2(n63), .B(n416), .Y(c[76]) );
  NOR3x1f_ASAP7_6t_L U682 ( .A(n62), .B(n125), .C(n417), .Y(n416) );
  OAI22xp5_ASAP7_6t_L U683 ( .A1(n418), .A2(n419), .B1(n420), .B2(n421), .Y(
        n63) );
  INVx1_ASAP7_6t_L U684 ( .A(n420), .Y(n419) );
  INVx1_ASAP7_6t_L U685 ( .A(n422), .Y(n62) );
  XOR2xp5r_ASAP7_6t_L U686 ( .A(n362), .B(n423), .Y(n422) );
  XOR2xp5r_ASAP7_6t_L U687 ( .A(n424), .B(n364), .Y(n423) );
  XOR2xp5r_ASAP7_6t_L U688 ( .A(n365), .B(n425), .Y(n364) );
  XOR2xp5r_ASAP7_6t_L U689 ( .A(n413), .B(n414), .Y(n425) );
  XOR2xp5r_ASAP7_6t_L U690 ( .A(n426), .B(n415), .Y(n414) );
  XOR2xp5r_ASAP7_6t_L U691 ( .A(n374), .B(n369), .Y(n415) );
  XOR2xp5r_ASAP7_6t_L U692 ( .A(n373), .B(n427), .Y(n369) );
  XOR2xp5r_ASAP7_6t_L U693 ( .A(n376), .B(n375), .Y(n427) );
  AOI21xp25_ASAP7_6t_L U694 ( .A1(n428), .A2(n429), .B(n430), .Y(n375) );
  NOR3x1f_ASAP7_6t_L U695 ( .A(n429), .B(n250), .C(n170), .Y(n430) );
  XOR2xp5r_ASAP7_6t_L U696 ( .A(n378), .B(n431), .Y(n376) );
  XOR2xp5r_ASAP7_6t_L U697 ( .A(n381), .B(n380), .Y(n431) );
  INVx1_ASAP7_6t_L U698 ( .A(n382), .Y(n380) );
  XOR2xp5r_ASAP7_6t_L U699 ( .A(n432), .B(n383), .Y(n382) );
  XOR2xp5r_ASAP7_6t_L U700 ( .A(n396), .B(n395), .Y(n383) );
  NOR2xp5_ASAP7_6t_L U701 ( .A(n285), .B(n159), .Y(n395) );
  XOR2xp5r_ASAP7_6t_L U702 ( .A(n393), .B(n394), .Y(n396) );
  NOR2xp5_ASAP7_6t_L U703 ( .A(n433), .B(n113), .Y(n394) );
  NOR2xp5_ASAP7_6t_L U704 ( .A(n392), .B(n117), .Y(n393) );
  AOI21xp25_ASAP7_6t_L U705 ( .A1(n434), .A2(n435), .B(n436), .Y(n432) );
  NOR3x1f_ASAP7_6t_L U706 ( .A(n434), .B(n146), .C(n280), .Y(n436) );
  XOR2xp5r_ASAP7_6t_L U707 ( .A(n387), .B(n388), .Y(n381) );
  NAND2xp5R_ASAP7_6t_L U708 ( .A(b[10]), .B(a[9]), .Y(n388) );
  XOR2xp5r_ASAP7_6t_L U709 ( .A(n437), .B(n390), .Y(n387) );
  NAND2xp5R_ASAP7_6t_L U710 ( .A(b[11]), .B(a[8]), .Y(n390) );
  INVx1_ASAP7_6t_L U711 ( .A(n389), .Y(n437) );
  NAND2xp5R_ASAP7_6t_L U712 ( .A(a[7]), .B(b[12]), .Y(n389) );
  AOI22xp25_ASAP7_6t_L U713 ( .A1(n438), .A2(n439), .B1(n440), .B2(n441), .Y(
        n378) );
  AO21x1_ASAP7_6t_L U714 ( .A1(n442), .A2(n443), .B(n444), .Y(n373) );
  NOR3x1f_ASAP7_6t_L U715 ( .A(n442), .B(n126), .C(n285), .Y(n444) );
  OAI22xp5_ASAP7_6t_L U716 ( .A1(n445), .A2(n446), .B1(n447), .B2(n448), .Y(
        n374) );
  AOI21xp25_ASAP7_6t_L U717 ( .A1(n449), .A2(n450), .B(n451), .Y(n426) );
  NOR3x1f_ASAP7_6t_L U718 ( .A(n450), .B(n212), .C(n195), .Y(n451) );
  XOR2xp5r_ASAP7_6t_L U719 ( .A(n409), .B(n410), .Y(n413) );
  OAI22xp5_ASAP7_6t_L U720 ( .A1(n452), .A2(n453), .B1(n454), .B2(n455), .Y(
        n410) );
  INVx1_ASAP7_6t_L U721 ( .A(n453), .Y(n454) );
  XOR2xp5r_ASAP7_6t_L U722 ( .A(n456), .B(n397), .Y(n409) );
  AOI21xp25_ASAP7_6t_L U723 ( .A1(n457), .A2(n458), .B(n459), .Y(n397) );
  NOR3x1f_ASAP7_6t_L U724 ( .A(n458), .B(n114), .C(n311), .Y(n459) );
  XOR2xp5r_ASAP7_6t_L U725 ( .A(n460), .B(n398), .Y(n456) );
  XOR2xp5r_ASAP7_6t_L U726 ( .A(n461), .B(n403), .Y(n398) );
  XOR2xp5r_ASAP7_6t_L U727 ( .A(n462), .B(n402), .Y(n403) );
  NOR2xp5_ASAP7_6t_L U728 ( .A(n195), .B(n185), .Y(n402) );
  NAND2xp5R_ASAP7_6t_L U729 ( .A(a[11]), .B(b[8]), .Y(n462) );
  XOR2xp5r_ASAP7_6t_L U730 ( .A(n463), .B(n400), .Y(n461) );
  NAND2xp5R_ASAP7_6t_L U731 ( .A(b[6]), .B(a[13]), .Y(n400) );
  NAND2xp5R_ASAP7_6t_L U732 ( .A(b[7]), .B(a[12]), .Y(n463) );
  NOR2xp5_ASAP7_6t_L U733 ( .A(n131), .B(n361), .Y(n460) );
  AOI21xp25_ASAP7_6t_L U734 ( .A1(n464), .A2(n465), .B(n466), .Y(n365) );
  NOR3x1f_ASAP7_6t_L U735 ( .A(n464), .B(n131), .C(n417), .Y(n466) );
  NOR2xp5_ASAP7_6t_L U736 ( .A(n125), .B(n417), .Y(n424) );
  AOI22xp25_ASAP7_6t_L U737 ( .A1(n467), .A2(n468), .B1(n469), .B2(n470), .Y(
        n362) );
  AO21x1_ASAP7_6t_L U738 ( .A1(n64), .A2(n65), .B(n471), .Y(c[75]) );
  NOR3x1f_ASAP7_6t_L U739 ( .A(n65), .B(n125), .C(n472), .Y(n471) );
  XOR2xp5r_ASAP7_6t_L U740 ( .A(n421), .B(n473), .Y(n65) );
  XOR2xp5r_ASAP7_6t_L U741 ( .A(n474), .B(n420), .Y(n473) );
  XOR2xp5r_ASAP7_6t_L U742 ( .A(n418), .B(n475), .Y(n420) );
  XOR2xp5r_ASAP7_6t_L U743 ( .A(n468), .B(n467), .Y(n475) );
  INVx1_ASAP7_6t_L U744 ( .A(n470), .Y(n467) );
  XOR2xp5r_ASAP7_6t_L U745 ( .A(n476), .B(n469), .Y(n470) );
  XOR2xp5r_ASAP7_6t_L U746 ( .A(n450), .B(n449), .Y(n469) );
  OAI22xp5_ASAP7_6t_L U747 ( .A1(n477), .A2(n478), .B1(n479), .B2(n480), .Y(
        n449) );
  INVx1_ASAP7_6t_L U748 ( .A(n479), .Y(n478) );
  XOR2xp5r_ASAP7_6t_L U749 ( .A(n448), .B(n481), .Y(n450) );
  XOR2xp5r_ASAP7_6t_L U750 ( .A(n482), .B(n447), .Y(n481) );
  INVx1_ASAP7_6t_L U751 ( .A(n446), .Y(n447) );
  XOR2xp5r_ASAP7_6t_L U752 ( .A(n483), .B(n429), .Y(n446) );
  XOR2xp5r_ASAP7_6t_L U753 ( .A(n484), .B(n428), .Y(n429) );
  XOR2xp5r_ASAP7_6t_L U754 ( .A(n434), .B(n435), .Y(n428) );
  AO21x1_ASAP7_6t_L U755 ( .A1(n485), .A2(n486), .B(n487), .Y(n435) );
  NOR3x1f_ASAP7_6t_L U756 ( .A(n485), .B(n126), .C(n392), .Y(n487) );
  XOR2xp5r_ASAP7_6t_L U757 ( .A(n488), .B(n443), .Y(n434) );
  OAI22xp5_ASAP7_6t_L U758 ( .A1(n489), .A2(n490), .B1(n491), .B2(n492), .Y(
        n443) );
  XOR2xp5r_ASAP7_6t_L U759 ( .A(n493), .B(n442), .Y(n488) );
  XOR2xp5r_ASAP7_6t_L U760 ( .A(n438), .B(n494), .Y(n442) );
  XOR2xp5r_ASAP7_6t_L U761 ( .A(n495), .B(n439), .Y(n494) );
  NOR2xp5_ASAP7_6t_L U762 ( .A(n392), .B(n159), .Y(n439) );
  NOR2xp5_ASAP7_6t_L U763 ( .A(n126), .B(n285), .Y(n495) );
  INVx1_ASAP7_6t_L U764 ( .A(n440), .Y(n438) );
  XOR2xp5r_ASAP7_6t_L U765 ( .A(n441), .B(n496), .Y(n440) );
  NAND2xp5R_ASAP7_6t_L U766 ( .A(a[4]), .B(b[14]), .Y(n496) );
  NOR2xp5_ASAP7_6t_L U767 ( .A(n497), .B(n113), .Y(n441) );
  NOR2xp5_ASAP7_6t_L U768 ( .A(n146), .B(n280), .Y(n493) );
  AOI21xp25_ASAP7_6t_L U769 ( .A1(n498), .A2(n499), .B(n500), .Y(n484) );
  NOR3x1f_ASAP7_6t_L U770 ( .A(n498), .B(n146), .C(n285), .Y(n500) );
  XOR2xp5r_ASAP7_6t_L U771 ( .A(n445), .B(n501), .Y(n483) );
  NOR2xp5_ASAP7_6t_L U772 ( .A(n250), .B(n170), .Y(n501) );
  AOI22xp25_ASAP7_6t_L U773 ( .A1(n502), .A2(n503), .B1(n504), .B2(n505), .Y(
        n445) );
  NOR2xp5_ASAP7_6t_L U774 ( .A(n212), .B(n195), .Y(n482) );
  AOI22xp25_ASAP7_6t_L U775 ( .A1(n506), .A2(n507), .B1(n508), .B2(n509), .Y(
        n448) );
  AOI21xp25_ASAP7_6t_L U776 ( .A1(n510), .A2(n511), .B(n512), .Y(n476) );
  NOR3x1f_ASAP7_6t_L U777 ( .A(n511), .B(n185), .C(n296), .Y(n512) );
  XOR2xp5r_ASAP7_6t_L U778 ( .A(n464), .B(n465), .Y(n468) );
  OAI22xp5_ASAP7_6t_L U779 ( .A1(n513), .A2(n514), .B1(n515), .B2(n516), .Y(
        n465) );
  INVx1_ASAP7_6t_L U780 ( .A(n514), .Y(n515) );
  XOR2xp5r_ASAP7_6t_L U781 ( .A(n517), .B(n452), .Y(n464) );
  AOI21xp25_ASAP7_6t_L U782 ( .A1(n518), .A2(n519), .B(n520), .Y(n452) );
  NOR3x1f_ASAP7_6t_L U783 ( .A(n519), .B(n114), .C(n361), .Y(n520) );
  XOR2xp5r_ASAP7_6t_L U784 ( .A(n521), .B(n453), .Y(n517) );
  XOR2xp5r_ASAP7_6t_L U785 ( .A(n458), .B(n522), .Y(n453) );
  XOR2xp5r_ASAP7_6t_L U786 ( .A(n455), .B(n523), .Y(n522) );
  NAND2xp5R_ASAP7_6t_L U787 ( .A(b[6]), .B(a[12]), .Y(n523) );
  NAND2xp5R_ASAP7_6t_L U788 ( .A(b[5]), .B(a[13]), .Y(n455) );
  XOR2xp5r_ASAP7_6t_L U789 ( .A(n524), .B(n457), .Y(n458) );
  NOR2xp5_ASAP7_6t_L U790 ( .A(n258), .B(n185), .Y(n457) );
  NAND2xp5R_ASAP7_6t_L U791 ( .A(a[11]), .B(b[7]), .Y(n524) );
  NOR2xp5_ASAP7_6t_L U792 ( .A(n131), .B(n417), .Y(n521) );
  AOI21xp25_ASAP7_6t_L U793 ( .A1(n525), .A2(n526), .B(n527), .Y(n418) );
  NOR3x1f_ASAP7_6t_L U794 ( .A(n525), .B(n131), .C(n472), .Y(n527) );
  NOR2xp5_ASAP7_6t_L U795 ( .A(n125), .B(n472), .Y(n474) );
  AOI22xp25_ASAP7_6t_L U796 ( .A1(n528), .A2(n529), .B1(n530), .B2(n531), .Y(
        n421) );
  INVx1_ASAP7_6t_L U797 ( .A(n530), .Y(n529) );
  OAI22xp5_ASAP7_6t_L U798 ( .A1(n532), .A2(n533), .B1(n534), .B2(n535), .Y(
        n64) );
  INVx1_ASAP7_6t_L U799 ( .A(n533), .Y(n534) );
  AO21x1_ASAP7_6t_L U800 ( .A1(n67), .A2(n66), .B(n536), .Y(c[74]) );
  NOR3x1f_ASAP7_6t_L U801 ( .A(n67), .B(n125), .C(n537), .Y(n536) );
  OAI22xp5_ASAP7_6t_L U802 ( .A1(n538), .A2(n539), .B1(n540), .B2(n541), .Y(
        n66) );
  INVx1_ASAP7_6t_L U803 ( .A(n539), .Y(n540) );
  XOR2xp5r_ASAP7_6t_L U804 ( .A(n532), .B(n542), .Y(n67) );
  XOR2xp5r_ASAP7_6t_L U805 ( .A(n543), .B(n533), .Y(n542) );
  XOR2xp5r_ASAP7_6t_L U806 ( .A(n535), .B(n544), .Y(n533) );
  XOR2xp5r_ASAP7_6t_L U807 ( .A(n531), .B(n530), .Y(n544) );
  OAI22xp5_ASAP7_6t_L U808 ( .A1(n545), .A2(n546), .B1(n547), .B2(n548), .Y(
        n530) );
  XOR2xp5r_ASAP7_6t_L U809 ( .A(n549), .B(n550), .Y(n548) );
  INVx1_ASAP7_6t_L U810 ( .A(n546), .Y(n547) );
  XOR2xp5r_ASAP7_6t_L U811 ( .A(n551), .B(n550), .Y(n545) );
  INVx1_ASAP7_6t_L U812 ( .A(n528), .Y(n550) );
  XOR2xp5r_ASAP7_6t_L U813 ( .A(n510), .B(n511), .Y(n528) );
  XOR2xp5r_ASAP7_6t_L U814 ( .A(n480), .B(n552), .Y(n511) );
  XOR2xp5r_ASAP7_6t_L U815 ( .A(n553), .B(n479), .Y(n552) );
  XOR2xp5r_ASAP7_6t_L U816 ( .A(n507), .B(n554), .Y(n479) );
  XOR2xp5r_ASAP7_6t_L U817 ( .A(n477), .B(n506), .Y(n554) );
  INVx1_ASAP7_6t_L U818 ( .A(n508), .Y(n506) );
  XOR2xp5r_ASAP7_6t_L U819 ( .A(n555), .B(n509), .Y(n508) );
  XOR2xp5r_ASAP7_6t_L U820 ( .A(n499), .B(n498), .Y(n509) );
  XOR2xp5r_ASAP7_6t_L U821 ( .A(n556), .B(n486), .Y(n498) );
  AO21x1_ASAP7_6t_L U822 ( .A1(n557), .A2(n558), .B(n559), .Y(n486) );
  NOR3x1f_ASAP7_6t_L U823 ( .A(n558), .B(n159), .C(n497), .Y(n559) );
  XOR2xp5r_ASAP7_6t_L U824 ( .A(n560), .B(n485), .Y(n556) );
  XOR2xp5r_ASAP7_6t_L U825 ( .A(n561), .B(n491), .Y(n485) );
  INVx1_ASAP7_6t_L U826 ( .A(n489), .Y(n491) );
  XOR2xp5r_ASAP7_6t_L U827 ( .A(n562), .B(n492), .Y(n489) );
  NAND2xp5R_ASAP7_6t_L U828 ( .A(a[2]), .B(b[15]), .Y(n492) );
  NOR2xp5_ASAP7_6t_L U829 ( .A(n117), .B(n497), .Y(n562) );
  XOR2xp5r_ASAP7_6t_L U830 ( .A(n563), .B(n490), .Y(n561) );
  NAND2xp5R_ASAP7_6t_L U831 ( .A(a[4]), .B(b[13]), .Y(n490) );
  NAND2xp5R_ASAP7_6t_L U832 ( .A(a[5]), .B(b[12]), .Y(n563) );
  NOR2xp5_ASAP7_6t_L U833 ( .A(n146), .B(n285), .Y(n560) );
  OAI22xp5_ASAP7_6t_L U834 ( .A1(n564), .A2(n565), .B1(n566), .B2(n567), .Y(
        n499) );
  AOI21xp25_ASAP7_6t_L U835 ( .A1(n568), .A2(n569), .B(n570), .Y(n555) );
  NOR3x1f_ASAP7_6t_L U836 ( .A(n568), .B(n146), .C(n392), .Y(n570) );
  AOI22xp25_ASAP7_6t_L U837 ( .A1(n571), .A2(n572), .B1(n573), .B2(n574), .Y(
        n477) );
  XOR2xp5r_ASAP7_6t_L U838 ( .A(n502), .B(n503), .Y(n507) );
  NOR2xp5_ASAP7_6t_L U839 ( .A(n258), .B(n212), .Y(n503) );
  XOR2xp5r_ASAP7_6t_L U840 ( .A(n505), .B(n504), .Y(n502) );
  NOR2xp5_ASAP7_6t_L U841 ( .A(n170), .B(n280), .Y(n504) );
  NOR2xp5_ASAP7_6t_L U842 ( .A(n195), .B(n250), .Y(n505) );
  NOR2xp5_ASAP7_6t_L U843 ( .A(n185), .B(n296), .Y(n553) );
  AOI22xp25_ASAP7_6t_L U844 ( .A1(n575), .A2(n576), .B1(n577), .B2(n578), .Y(
        n480) );
  OAI22xp5_ASAP7_6t_L U845 ( .A1(n579), .A2(n580), .B1(n581), .B2(n582), .Y(
        n510) );
  INVx1_ASAP7_6t_L U846 ( .A(n581), .Y(n580) );
  XOR2xp5r_ASAP7_6t_L U847 ( .A(n526), .B(n525), .Y(n531) );
  XOR2xp5r_ASAP7_6t_L U848 ( .A(n513), .B(n583), .Y(n525) );
  XOR2xp5r_ASAP7_6t_L U849 ( .A(n584), .B(n514), .Y(n583) );
  XOR2xp5r_ASAP7_6t_L U850 ( .A(n585), .B(n519), .Y(n514) );
  XOR2xp5r_ASAP7_6t_L U851 ( .A(n518), .B(n586), .Y(n519) );
  NAND2xp5R_ASAP7_6t_L U852 ( .A(b[6]), .B(a[11]), .Y(n586) );
  NOR3x1f_ASAP7_6t_L U853 ( .A(n587), .B(n185), .C(n311), .Y(n518) );
  XOR2xp5r_ASAP7_6t_L U854 ( .A(n588), .B(n516), .Y(n585) );
  NAND2xp5R_ASAP7_6t_L U855 ( .A(b[4]), .B(a[13]), .Y(n516) );
  NAND2xp5R_ASAP7_6t_L U856 ( .A(b[5]), .B(a[12]), .Y(n588) );
  NOR2xp5_ASAP7_6t_L U857 ( .A(n131), .B(n472), .Y(n584) );
  AOI21xp25_ASAP7_6t_L U858 ( .A1(n589), .A2(n590), .B(n591), .Y(n513) );
  NOR3x1f_ASAP7_6t_L U859 ( .A(n590), .B(n114), .C(n417), .Y(n591) );
  OAI22xp5_ASAP7_6t_L U860 ( .A1(n592), .A2(n593), .B1(n594), .B2(n595), .Y(
        n526) );
  INVx1_ASAP7_6t_L U861 ( .A(n593), .Y(n594) );
  AOI21xp25_ASAP7_6t_L U862 ( .A1(n596), .A2(n597), .B(n598), .Y(n535) );
  NOR3x1f_ASAP7_6t_L U863 ( .A(n596), .B(n131), .C(n537), .Y(n598) );
  NOR2xp5_ASAP7_6t_L U864 ( .A(n125), .B(n537), .Y(n543) );
  AOI22xp25_ASAP7_6t_L U865 ( .A1(n599), .A2(n600), .B1(n601), .B2(n602), .Y(
        n532) );
  INVx1_ASAP7_6t_L U866 ( .A(n601), .Y(n600) );
  AO21x1_ASAP7_6t_L U867 ( .A1(n69), .A2(n68), .B(n603), .Y(c[73]) );
  NOR3x1f_ASAP7_6t_L U868 ( .A(n69), .B(n125), .C(n99), .Y(n603) );
  OAI22xp5_ASAP7_6t_L U869 ( .A1(n604), .A2(n605), .B1(n606), .B2(n607), .Y(
        n68) );
  INVx1_ASAP7_6t_L U870 ( .A(n606), .Y(n605) );
  XOR2xp5r_ASAP7_6t_L U871 ( .A(n538), .B(n608), .Y(n69) );
  XOR2xp5r_ASAP7_6t_L U872 ( .A(n609), .B(n539), .Y(n608) );
  XOR2xp5r_ASAP7_6t_L U873 ( .A(n541), .B(n610), .Y(n539) );
  XOR2xp5r_ASAP7_6t_L U874 ( .A(n602), .B(n601), .Y(n610) );
  OAI22xp5_ASAP7_6t_L U875 ( .A1(n611), .A2(n612), .B1(n613), .B2(n614), .Y(
        n601) );
  XOR2xp5r_ASAP7_6t_L U876 ( .A(n615), .B(n599), .Y(n614) );
  XOR2xp5r_ASAP7_6t_L U877 ( .A(n616), .B(n599), .Y(n611) );
  XOR2xp5r_ASAP7_6t_L U878 ( .A(n549), .B(n546), .Y(n599) );
  XOR2xp5r_ASAP7_6t_L U879 ( .A(n582), .B(n617), .Y(n546) );
  XOR2xp5r_ASAP7_6t_L U880 ( .A(n551), .B(n581), .Y(n617) );
  XOR2xp5r_ASAP7_6t_L U881 ( .A(n576), .B(n618), .Y(n581) );
  XOR2xp5r_ASAP7_6t_L U882 ( .A(n579), .B(n575), .Y(n618) );
  INVx1_ASAP7_6t_L U883 ( .A(n577), .Y(n575) );
  XOR2xp5r_ASAP7_6t_L U884 ( .A(n619), .B(n578), .Y(n577) );
  XOR2xp5r_ASAP7_6t_L U885 ( .A(n568), .B(n569), .Y(n578) );
  OAI22xp5_ASAP7_6t_L U886 ( .A1(n620), .A2(n621), .B1(n622), .B2(n623), .Y(
        n569) );
  INVx1_ASAP7_6t_L U887 ( .A(n621), .Y(n622) );
  XOR2xp5r_ASAP7_6t_L U888 ( .A(n624), .B(n564), .Y(n568) );
  AOI21xp25_ASAP7_6t_L U889 ( .A1(n625), .A2(n626), .B(n627), .Y(n564) );
  NOR3x1f_ASAP7_6t_L U890 ( .A(n626), .B(n159), .C(n96), .Y(n627) );
  XOR2xp5r_ASAP7_6t_L U891 ( .A(n628), .B(n565), .Y(n624) );
  INVx1_ASAP7_6t_L U892 ( .A(n566), .Y(n565) );
  XOR2xp5r_ASAP7_6t_L U893 ( .A(n558), .B(n629), .Y(n566) );
  XOR2xp5r_ASAP7_6t_L U894 ( .A(n630), .B(n567), .Y(n629) );
  NAND2xp5R_ASAP7_6t_L U895 ( .A(a[4]), .B(b[12]), .Y(n567) );
  NOR2xp5_ASAP7_6t_L U896 ( .A(n159), .B(n497), .Y(n630) );
  XOR2xp5r_ASAP7_6t_L U897 ( .A(n557), .B(n631), .Y(n558) );
  NAND2xp5R_ASAP7_6t_L U898 ( .A(a[2]), .B(b[14]), .Y(n631) );
  NOR2xp5_ASAP7_6t_L U899 ( .A(n100), .B(n113), .Y(n557) );
  NOR2xp5_ASAP7_6t_L U900 ( .A(n146), .B(n392), .Y(n628) );
  AOI21xp25_ASAP7_6t_L U901 ( .A1(n632), .A2(n633), .B(n634), .Y(n619) );
  NOR3x1f_ASAP7_6t_L U902 ( .A(n632), .B(n146), .C(n433), .Y(n634) );
  AOI22xp25_ASAP7_6t_L U903 ( .A1(n635), .A2(n636), .B1(n637), .B2(n638), .Y(
        n579) );
  XOR2xp5r_ASAP7_6t_L U904 ( .A(n571), .B(n572), .Y(n576) );
  NOR2xp5_ASAP7_6t_L U905 ( .A(n258), .B(n250), .Y(n572) );
  XOR2xp5r_ASAP7_6t_L U906 ( .A(n574), .B(n573), .Y(n571) );
  NOR2xp5_ASAP7_6t_L U907 ( .A(n170), .B(n285), .Y(n573) );
  NOR2xp5_ASAP7_6t_L U908 ( .A(n195), .B(n280), .Y(n574) );
  XOR2xp5r_ASAP7_6t_L U909 ( .A(n639), .B(n587), .Y(n551) );
  NAND2xp5R_ASAP7_6t_L U910 ( .A(b[7]), .B(a[9]), .Y(n587) );
  NAND2xp5R_ASAP7_6t_L U911 ( .A(a[10]), .B(b[6]), .Y(n639) );
  AOI22xp25_ASAP7_6t_L U912 ( .A1(n640), .A2(n641), .B1(n642), .B2(n643), .Y(
        n582) );
  OAI22xp5_ASAP7_6t_L U913 ( .A1(n644), .A2(n645), .B1(n646), .B2(n647), .Y(
        n549) );
  XOR2xp5r_ASAP7_6t_L U914 ( .A(n597), .B(n596), .Y(n602) );
  XOR2xp5r_ASAP7_6t_L U915 ( .A(n592), .B(n648), .Y(n596) );
  XOR2xp5r_ASAP7_6t_L U916 ( .A(n649), .B(n593), .Y(n648) );
  XOR2xp5r_ASAP7_6t_L U917 ( .A(n650), .B(n590), .Y(n593) );
  XOR2xp5r_ASAP7_6t_L U918 ( .A(n589), .B(n651), .Y(n590) );
  NAND2xp5R_ASAP7_6t_L U919 ( .A(b[5]), .B(a[11]), .Y(n651) );
  NOR3x1f_ASAP7_6t_L U920 ( .A(n652), .B(n212), .C(n311), .Y(n589) );
  XOR2xp5r_ASAP7_6t_L U921 ( .A(n653), .B(n595), .Y(n650) );
  NAND2xp5R_ASAP7_6t_L U922 ( .A(b[3]), .B(a[13]), .Y(n595) );
  NAND2xp5R_ASAP7_6t_L U923 ( .A(b[4]), .B(a[12]), .Y(n653) );
  NOR2xp5_ASAP7_6t_L U924 ( .A(n131), .B(n537), .Y(n649) );
  AOI21xp25_ASAP7_6t_L U925 ( .A1(n654), .A2(n655), .B(n656), .Y(n592) );
  NOR3x1f_ASAP7_6t_L U926 ( .A(n655), .B(n114), .C(n472), .Y(n656) );
  OAI22xp5_ASAP7_6t_L U927 ( .A1(n657), .A2(n658), .B1(n659), .B2(n660), .Y(
        n597) );
  INVx1_ASAP7_6t_L U928 ( .A(n658), .Y(n659) );
  AOI21xp25_ASAP7_6t_L U929 ( .A1(n661), .A2(n662), .B(n663), .Y(n541) );
  NOR3x1f_ASAP7_6t_L U930 ( .A(n661), .B(n131), .C(n99), .Y(n663) );
  NOR2xp5_ASAP7_6t_L U931 ( .A(n125), .B(n99), .Y(n609) );
  AOI22xp25_ASAP7_6t_L U932 ( .A1(n664), .A2(n665), .B1(n666), .B2(n667), .Y(
        n538) );
  AO21x1_ASAP7_6t_L U933 ( .A1(n70), .A2(n71), .B(n668), .Y(c[72]) );
  NOR3x1f_ASAP7_6t_L U934 ( .A(n71), .B(n125), .C(n97), .Y(n668) );
  XOR2xp5r_ASAP7_6t_L U935 ( .A(n607), .B(n669), .Y(n71) );
  XOR2xp5r_ASAP7_6t_L U936 ( .A(n670), .B(n606), .Y(n669) );
  XOR2xp5r_ASAP7_6t_L U937 ( .A(n604), .B(n671), .Y(n606) );
  XOR2xp5r_ASAP7_6t_L U938 ( .A(n665), .B(n664), .Y(n671) );
  INVx1_ASAP7_6t_L U939 ( .A(n667), .Y(n664) );
  XOR2xp5r_ASAP7_6t_L U940 ( .A(n672), .B(n666), .Y(n667) );
  XOR2xp5r_ASAP7_6t_L U941 ( .A(n615), .B(n613), .Y(n666) );
  INVx1_ASAP7_6t_L U942 ( .A(n612), .Y(n613) );
  XOR2xp5r_ASAP7_6t_L U943 ( .A(n647), .B(n673), .Y(n612) );
  XOR2xp5r_ASAP7_6t_L U944 ( .A(n616), .B(n645), .Y(n673) );
  INVx1_ASAP7_6t_L U945 ( .A(n646), .Y(n645) );
  XOR2xp5r_ASAP7_6t_L U946 ( .A(n641), .B(n674), .Y(n646) );
  XOR2xp5r_ASAP7_6t_L U947 ( .A(n644), .B(n640), .Y(n674) );
  INVx1_ASAP7_6t_L U948 ( .A(n642), .Y(n640) );
  XOR2xp5r_ASAP7_6t_L U949 ( .A(n675), .B(n643), .Y(n642) );
  XOR2xp5r_ASAP7_6t_L U950 ( .A(n632), .B(n633), .Y(n643) );
  OAI22xp5_ASAP7_6t_L U951 ( .A1(n676), .A2(n677), .B1(n678), .B2(n679), .Y(
        n633) );
  XOR2xp5r_ASAP7_6t_L U952 ( .A(n680), .B(n620), .Y(n632) );
  AOI21xp25_ASAP7_6t_L U953 ( .A1(n681), .A2(n682), .B(n683), .Y(n620) );
  NOR3x1f_ASAP7_6t_L U954 ( .A(n682), .B(n126), .C(n96), .Y(n683) );
  XOR2xp5r_ASAP7_6t_L U955 ( .A(n684), .B(n621), .Y(n680) );
  XOR2xp5r_ASAP7_6t_L U956 ( .A(n685), .B(n626), .Y(n621) );
  XOR2xp5r_ASAP7_6t_L U957 ( .A(n686), .B(n625), .Y(n626) );
  NOR2xp5_ASAP7_6t_L U958 ( .A(n98), .B(n113), .Y(n625) );
  INVx1_ASAP7_6t_L U959 ( .A(b[15]), .Y(n113) );
  NAND2xp5R_ASAP7_6t_L U960 ( .A(b[14]), .B(a[1]), .Y(n686) );
  XOR2xp5r_ASAP7_6t_L U961 ( .A(n687), .B(n623), .Y(n685) );
  NAND2xp5R_ASAP7_6t_L U962 ( .A(a[3]), .B(b[12]), .Y(n623) );
  NAND2xp5R_ASAP7_6t_L U963 ( .A(a[2]), .B(b[13]), .Y(n687) );
  NOR2xp5_ASAP7_6t_L U964 ( .A(n146), .B(n433), .Y(n684) );
  NOR2xp5_ASAP7_6t_L U965 ( .A(n688), .B(n689), .Y(n675) );
  NOR3x1f_ASAP7_6t_L U966 ( .A(n690), .B(n691), .C(n692), .Y(n689) );
  NOR3x1f_ASAP7_6t_L U967 ( .A(n693), .B(n170), .C(n433), .Y(n688) );
  AOI22xp25_ASAP7_6t_L U968 ( .A1(n694), .A2(n695), .B1(n696), .B2(n697), .Y(
        n644) );
  XOR2xp5r_ASAP7_6t_L U969 ( .A(n635), .B(n636), .Y(n641) );
  NOR2xp5_ASAP7_6t_L U970 ( .A(n258), .B(n280), .Y(n636) );
  XOR2xp5r_ASAP7_6t_L U971 ( .A(n638), .B(n637), .Y(n635) );
  NOR2xp5_ASAP7_6t_L U972 ( .A(n170), .B(n392), .Y(n637) );
  NOR2xp5_ASAP7_6t_L U973 ( .A(n195), .B(n285), .Y(n638) );
  XOR2xp5r_ASAP7_6t_L U974 ( .A(n698), .B(n699), .Y(n616) );
  NAND2xp5R_ASAP7_6t_L U975 ( .A(b[6]), .B(a[9]), .Y(n699) );
  INVx1_ASAP7_6t_L U976 ( .A(n652), .Y(n698) );
  NAND2xp5R_ASAP7_6t_L U977 ( .A(b[7]), .B(a[8]), .Y(n652) );
  AOI22xp25_ASAP7_6t_L U978 ( .A1(n700), .A2(n701), .B1(n702), .B2(n703), .Y(
        n647) );
  INVx1_ASAP7_6t_L U979 ( .A(n700), .Y(n702) );
  AOI22xp25_ASAP7_6t_L U980 ( .A1(n704), .A2(n705), .B1(n706), .B2(n707), .Y(
        n615) );
  INVx1_ASAP7_6t_L U981 ( .A(n705), .Y(n706) );
  AOI21xp25_ASAP7_6t_L U982 ( .A1(n708), .A2(n709), .B(n710), .Y(n672) );
  NOR3x1f_ASAP7_6t_L U983 ( .A(n708), .B(n250), .C(n311), .Y(n710) );
  XOR2xp5r_ASAP7_6t_L U984 ( .A(n661), .B(n662), .Y(n665) );
  OAI22xp5_ASAP7_6t_L U985 ( .A1(n711), .A2(n712), .B1(n713), .B2(n714), .Y(
        n662) );
  XOR2xp5r_ASAP7_6t_L U986 ( .A(n715), .B(n657), .Y(n661) );
  AOI21xp25_ASAP7_6t_L U987 ( .A1(n716), .A2(n717), .B(n718), .Y(n657) );
  NOR3x1f_ASAP7_6t_L U988 ( .A(n717), .B(n160), .C(n472), .Y(n718) );
  XOR2xp5r_ASAP7_6t_L U989 ( .A(n719), .B(n658), .Y(n715) );
  XOR2xp5r_ASAP7_6t_L U990 ( .A(n720), .B(n655), .Y(n658) );
  XOR2xp5r_ASAP7_6t_L U991 ( .A(n721), .B(n654), .Y(n655) );
  NOR2xp5_ASAP7_6t_L U992 ( .A(n361), .B(n185), .Y(n654) );
  NAND2xp5R_ASAP7_6t_L U993 ( .A(a[11]), .B(b[4]), .Y(n721) );
  XOR2xp5r_ASAP7_6t_L U994 ( .A(n722), .B(n660), .Y(n720) );
  NAND2xp5R_ASAP7_6t_L U995 ( .A(b[2]), .B(a[13]), .Y(n660) );
  NAND2xp5R_ASAP7_6t_L U996 ( .A(b[3]), .B(a[12]), .Y(n722) );
  NOR2xp5_ASAP7_6t_L U997 ( .A(n131), .B(n99), .Y(n719) );
  AOI21xp25_ASAP7_6t_L U998 ( .A1(n723), .A2(n724), .B(n725), .Y(n604) );
  NOR3x1f_ASAP7_6t_L U999 ( .A(n723), .B(n116), .C(n99), .Y(n725) );
  NOR2xp5_ASAP7_6t_L U1000 ( .A(n125), .B(n97), .Y(n670) );
  INVx1_ASAP7_6t_L U1001 ( .A(a[15]), .Y(n125) );
  AOI22xp25_ASAP7_6t_L U1002 ( .A1(n726), .A2(n727), .B1(n728), .B2(n729), .Y(
        n607) );
  INVx1_ASAP7_6t_L U1003 ( .A(n728), .Y(n726) );
  OAI22xp5_ASAP7_6t_L U1004 ( .A1(n730), .A2(n731), .B1(n732), .B2(n733), .Y(
        n70) );
  INVx1_ASAP7_6t_L U1005 ( .A(n732), .Y(n731) );
  AO21x1_ASAP7_6t_L U1006 ( .A1(n73), .A2(n72), .B(n734), .Y(c[71]) );
  NOR3x1f_ASAP7_6t_L U1007 ( .A(n73), .B(n131), .C(n97), .Y(n734) );
  OAI22xp5_ASAP7_6t_L U1008 ( .A1(n735), .A2(n736), .B1(n737), .B2(n738), .Y(
        n72) );
  INVx1_ASAP7_6t_L U1009 ( .A(n736), .Y(n737) );
  XOR2xp5r_ASAP7_6t_L U1010 ( .A(n739), .B(n740), .Y(n73) );
  XOR2xp5r_ASAP7_6t_L U1011 ( .A(n741), .B(n732), .Y(n740) );
  XOR2xp5r_ASAP7_6t_L U1012 ( .A(n733), .B(n742), .Y(n732) );
  XOR2xp5r_ASAP7_6t_L U1013 ( .A(n727), .B(n728), .Y(n742) );
  XOR2xp5r_ASAP7_6t_L U1014 ( .A(n743), .B(n729), .Y(n728) );
  XOR2xp5r_ASAP7_6t_L U1015 ( .A(n709), .B(n708), .Y(n729) );
  XOR2xp5r_ASAP7_6t_L U1016 ( .A(n704), .B(n744), .Y(n708) );
  XOR2xp5r_ASAP7_6t_L U1017 ( .A(n745), .B(n705), .Y(n744) );
  XOR2xp5r_ASAP7_6t_L U1018 ( .A(n701), .B(n746), .Y(n705) );
  XOR2xp5r_ASAP7_6t_L U1019 ( .A(n707), .B(n700), .Y(n746) );
  XOR2xp5r_ASAP7_6t_L U1020 ( .A(n747), .B(n703), .Y(n700) );
  XOR2xp5r_ASAP7_6t_L U1021 ( .A(n748), .B(n693), .Y(n703) );
  INVx1_ASAP7_6t_L U1022 ( .A(n690), .Y(n693) );
  XOR2xp5r_ASAP7_6t_L U1023 ( .A(n749), .B(n676), .Y(n690) );
  AOI21xp25_ASAP7_6t_L U1024 ( .A1(n750), .A2(n751), .B(n752), .Y(n676) );
  NOR3x1f_ASAP7_6t_L U1025 ( .A(n751), .B(n146), .C(n96), .Y(n752) );
  XOR2xp5r_ASAP7_6t_L U1026 ( .A(n753), .B(n678), .Y(n749) );
  INVx1_ASAP7_6t_L U1027 ( .A(n677), .Y(n678) );
  XOR2xp5r_ASAP7_6t_L U1028 ( .A(n754), .B(n682), .Y(n677) );
  XOR2xp5r_ASAP7_6t_L U1029 ( .A(n681), .B(n755), .Y(n682) );
  NAND2xp5R_ASAP7_6t_L U1030 ( .A(a[1]), .B(b[13]), .Y(n755) );
  NOR2xp5_ASAP7_6t_L U1031 ( .A(n98), .B(n117), .Y(n681) );
  INVx1_ASAP7_6t_L U1032 ( .A(b[14]), .Y(n117) );
  XOR2xp5r_ASAP7_6t_L U1033 ( .A(n756), .B(n679), .Y(n754) );
  NAND2xp5R_ASAP7_6t_L U1034 ( .A(a[3]), .B(b[11]), .Y(n679) );
  NAND2xp5R_ASAP7_6t_L U1035 ( .A(a[2]), .B(b[12]), .Y(n756) );
  NOR2xp5_ASAP7_6t_L U1036 ( .A(n170), .B(n433), .Y(n753) );
  NOR2xp5_ASAP7_6t_L U1037 ( .A(n692), .B(n691), .Y(n748) );
  INVx1_ASAP7_6t_L U1038 ( .A(n757), .Y(n691) );
  NOR2xp5_ASAP7_6t_L U1039 ( .A(n758), .B(n759), .Y(n747) );
  NOR3x1f_ASAP7_6t_L U1040 ( .A(n760), .B(n285), .C(n296), .Y(n707) );
  XOR2xp5r_ASAP7_6t_L U1041 ( .A(n694), .B(n695), .Y(n701) );
  NOR2xp5_ASAP7_6t_L U1042 ( .A(n296), .B(n280), .Y(n695) );
  XOR2xp5r_ASAP7_6t_L U1043 ( .A(n697), .B(n696), .Y(n694) );
  NOR2xp5_ASAP7_6t_L U1044 ( .A(n195), .B(n392), .Y(n696) );
  NOR2xp5_ASAP7_6t_L U1045 ( .A(n258), .B(n285), .Y(n697) );
  NOR2xp5_ASAP7_6t_L U1046 ( .A(n250), .B(n311), .Y(n745) );
  OAI22xp5_ASAP7_6t_L U1047 ( .A1(n761), .A2(n762), .B1(n763), .B2(n764), .Y(
        n704) );
  INVx1_ASAP7_6t_L U1048 ( .A(n759), .Y(n762) );
  AO22x1_ASAP7_6t_L U1049 ( .A1(n765), .A2(n766), .B1(n767), .B2(n768), .Y(
        n709) );
  AOI21xp25_ASAP7_6t_L U1050 ( .A1(n769), .A2(n770), .B(n771), .Y(n743) );
  NOR3x1f_ASAP7_6t_L U1051 ( .A(n770), .B(n280), .C(n311), .Y(n771) );
  XOR2xp5r_ASAP7_6t_L U1052 ( .A(n724), .B(n723), .Y(n727) );
  XOR2xp5r_ASAP7_6t_L U1053 ( .A(n772), .B(n711), .Y(n723) );
  AOI21xp25_ASAP7_6t_L U1054 ( .A1(n773), .A2(n774), .B(n775), .Y(n711) );
  NOR3x1f_ASAP7_6t_L U1055 ( .A(n774), .B(n185), .C(n472), .Y(n775) );
  XOR2xp5r_ASAP7_6t_L U1056 ( .A(n776), .B(n712), .Y(n772) );
  INVx1_ASAP7_6t_L U1057 ( .A(n713), .Y(n712) );
  XOR2xp5r_ASAP7_6t_L U1058 ( .A(n717), .B(n777), .Y(n713) );
  XOR2xp5r_ASAP7_6t_L U1059 ( .A(n778), .B(n714), .Y(n777) );
  NAND2xp5R_ASAP7_6t_L U1060 ( .A(b[2]), .B(a[12]), .Y(n714) );
  NOR2xp5_ASAP7_6t_L U1061 ( .A(n160), .B(n472), .Y(n778) );
  XOR2xp5r_ASAP7_6t_L U1062 ( .A(n779), .B(n716), .Y(n717) );
  NOR2xp5_ASAP7_6t_L U1063 ( .A(n361), .B(n212), .Y(n716) );
  NAND2xp5R_ASAP7_6t_L U1064 ( .A(a[10]), .B(b[4]), .Y(n779) );
  NOR2xp5_ASAP7_6t_L U1065 ( .A(n116), .B(n99), .Y(n776) );
  OAI22xp5_ASAP7_6t_L U1066 ( .A1(n780), .A2(n781), .B1(n782), .B2(n783), .Y(
        n724) );
  AOI21xp25_ASAP7_6t_L U1067 ( .A1(n784), .A2(n785), .B(n786), .Y(n733) );
  NOR3x1f_ASAP7_6t_L U1068 ( .A(n784), .B(n114), .C(n99), .Y(n786) );
  NOR2xp5_ASAP7_6t_L U1069 ( .A(n131), .B(n97), .Y(n741) );
  INVx1_ASAP7_6t_L U1070 ( .A(a[14]), .Y(n131) );
  INVx1_ASAP7_6t_L U1071 ( .A(n730), .Y(n739) );
  AOI22xp25_ASAP7_6t_L U1072 ( .A1(n787), .A2(n788), .B1(n789), .B2(n790), .Y(
        n730) );
  INVx1_ASAP7_6t_L U1073 ( .A(n788), .Y(n789) );
  AO21x1_ASAP7_6t_L U1074 ( .A1(n74), .A2(n75), .B(n791), .Y(c[70]) );
  NOR3x1f_ASAP7_6t_L U1075 ( .A(n75), .B(n116), .C(n97), .Y(n791) );
  XOR2xp5r_ASAP7_6t_L U1076 ( .A(n792), .B(n793), .Y(n75) );
  XOR2xp5r_ASAP7_6t_L U1077 ( .A(n794), .B(n736), .Y(n793) );
  XOR2xp5r_ASAP7_6t_L U1078 ( .A(n735), .B(n795), .Y(n736) );
  XOR2xp5r_ASAP7_6t_L U1079 ( .A(n790), .B(n788), .Y(n795) );
  XOR2xp5r_ASAP7_6t_L U1080 ( .A(n796), .B(n787), .Y(n788) );
  XOR2xp5r_ASAP7_6t_L U1081 ( .A(n770), .B(n769), .Y(n787) );
  OAI21xp25_ASAP7_6t_L U1082 ( .A1(n797), .A2(n798), .B(n799), .Y(n769) );
  NAND3xp33R_ASAP7_6t_L U1083 ( .A(n797), .B(a[5]), .C(b[7]), .Y(n799) );
  XOR2xp5r_ASAP7_6t_L U1084 ( .A(n768), .B(n800), .Y(n770) );
  XOR2xp5r_ASAP7_6t_L U1085 ( .A(n801), .B(n767), .Y(n800) );
  INVx1_ASAP7_6t_L U1086 ( .A(n765), .Y(n767) );
  XOR2xp5r_ASAP7_6t_L U1087 ( .A(n764), .B(n802), .Y(n765) );
  XOR2xp5r_ASAP7_6t_L U1088 ( .A(n766), .B(n761), .Y(n802) );
  INVx1_ASAP7_6t_L U1089 ( .A(n763), .Y(n761) );
  XOR2xp5r_ASAP7_6t_L U1090 ( .A(n803), .B(n759), .Y(n763) );
  XOR2xp5r_ASAP7_6t_L U1091 ( .A(n757), .B(n758), .Y(n759) );
  NAND2xp5R_ASAP7_6t_L U1092 ( .A(a[4]), .B(b[9]), .Y(n758) );
  XOR2xp5r_ASAP7_6t_L U1093 ( .A(n751), .B(n804), .Y(n757) );
  XOR2xp5r_ASAP7_6t_L U1094 ( .A(n692), .B(n805), .Y(n804) );
  NAND2xp5R_ASAP7_6t_L U1095 ( .A(a[2]), .B(b[11]), .Y(n805) );
  NAND2xp5R_ASAP7_6t_L U1096 ( .A(a[3]), .B(b[10]), .Y(n692) );
  XOR2xp5r_ASAP7_6t_L U1097 ( .A(n806), .B(n750), .Y(n751) );
  NOR2xp5_ASAP7_6t_L U1098 ( .A(n98), .B(n159), .Y(n750) );
  INVx1_ASAP7_6t_L U1099 ( .A(b[13]), .Y(n159) );
  NAND2xp5R_ASAP7_6t_L U1100 ( .A(b[12]), .B(a[1]), .Y(n806) );
  AOI22xp25_ASAP7_6t_L U1101 ( .A1(n807), .A2(n808), .B1(n809), .B2(n810), .Y(
        n803) );
  NOR3x1f_ASAP7_6t_L U1102 ( .A(n811), .B(n258), .C(n433), .Y(n766) );
  XOR2xp5r_ASAP7_6t_L U1103 ( .A(n812), .B(n760), .Y(n764) );
  NAND2xp5R_ASAP7_6t_L U1104 ( .A(b[8]), .B(a[5]), .Y(n760) );
  NOR2xp5_ASAP7_6t_L U1105 ( .A(n285), .B(n296), .Y(n812) );
  NOR2xp5_ASAP7_6t_L U1106 ( .A(n280), .B(n311), .Y(n801) );
  AO22x1_ASAP7_6t_L U1107 ( .A1(n813), .A2(n814), .B1(n815), .B2(n816), .Y(
        n768) );
  AOI21xp25_ASAP7_6t_L U1108 ( .A1(n817), .A2(n818), .B(n819), .Y(n796) );
  NOR3x1f_ASAP7_6t_L U1109 ( .A(n817), .B(n285), .C(n311), .Y(n819) );
  XOR2xp5r_ASAP7_6t_L U1110 ( .A(n784), .B(n785), .Y(n790) );
  OAI22xp5_ASAP7_6t_L U1111 ( .A1(n820), .A2(n821), .B1(n822), .B2(n823), .Y(
        n785) );
  INVx1_ASAP7_6t_L U1112 ( .A(n821), .Y(n822) );
  XOR2xp5r_ASAP7_6t_L U1113 ( .A(n824), .B(n780), .Y(n784) );
  AOI21xp25_ASAP7_6t_L U1114 ( .A1(n825), .A2(n826), .B(n827), .Y(n780) );
  NOR3x1f_ASAP7_6t_L U1115 ( .A(n826), .B(n212), .C(n472), .Y(n827) );
  XOR2xp5r_ASAP7_6t_L U1116 ( .A(n828), .B(n781), .Y(n824) );
  INVx1_ASAP7_6t_L U1117 ( .A(n782), .Y(n781) );
  XOR2xp5r_ASAP7_6t_L U1118 ( .A(n774), .B(n829), .Y(n782) );
  XOR2xp5r_ASAP7_6t_L U1119 ( .A(n830), .B(n783), .Y(n829) );
  NAND2xp5R_ASAP7_6t_L U1120 ( .A(b[2]), .B(a[11]), .Y(n783) );
  NOR2xp5_ASAP7_6t_L U1121 ( .A(n185), .B(n472), .Y(n830) );
  XOR2xp5r_ASAP7_6t_L U1122 ( .A(n773), .B(n831), .Y(n774) );
  NAND2xp5R_ASAP7_6t_L U1123 ( .A(b[4]), .B(a[9]), .Y(n831) );
  NOR2xp5_ASAP7_6t_L U1124 ( .A(n361), .B(n250), .Y(n773) );
  NOR2xp5_ASAP7_6t_L U1125 ( .A(n114), .B(n99), .Y(n828) );
  AOI21xp25_ASAP7_6t_L U1126 ( .A1(n832), .A2(n833), .B(n834), .Y(n735) );
  NOR3x1f_ASAP7_6t_L U1127 ( .A(n832), .B(n160), .C(n99), .Y(n834) );
  NOR2xp5_ASAP7_6t_L U1128 ( .A(n116), .B(n97), .Y(n794) );
  INVx1_ASAP7_6t_L U1129 ( .A(a[13]), .Y(n116) );
  INVx1_ASAP7_6t_L U1130 ( .A(n738), .Y(n792) );
  AOI22xp25_ASAP7_6t_L U1131 ( .A1(n835), .A2(n836), .B1(n837), .B2(n838), .Y(
        n738) );
  OAI22xp5_ASAP7_6t_L U1132 ( .A1(n839), .A2(n840), .B1(n841), .B2(n842), .Y(
        n74) );
  INVx1_ASAP7_6t_L U1133 ( .A(n840), .Y(n841) );
  AO21x1_ASAP7_6t_L U1134 ( .A1(n77), .A2(n76), .B(n843), .Y(c[69]) );
  NOR3x1f_ASAP7_6t_L U1135 ( .A(n77), .B(n114), .C(n97), .Y(n843) );
  OAI22xp5_ASAP7_6t_L U1136 ( .A1(n844), .A2(n845), .B1(n846), .B2(n847), .Y(
        n76) );
  INVx1_ASAP7_6t_L U1137 ( .A(n845), .Y(n846) );
  XOR2xp5r_ASAP7_6t_L U1138 ( .A(n839), .B(n848), .Y(n77) );
  XOR2xp5r_ASAP7_6t_L U1139 ( .A(n849), .B(n840), .Y(n848) );
  XOR2xp5r_ASAP7_6t_L U1140 ( .A(n842), .B(n850), .Y(n840) );
  XOR2xp5r_ASAP7_6t_L U1141 ( .A(n836), .B(n835), .Y(n850) );
  INVx1_ASAP7_6t_L U1142 ( .A(n837), .Y(n835) );
  XOR2xp5r_ASAP7_6t_L U1143 ( .A(n851), .B(n838), .Y(n837) );
  XOR2xp5r_ASAP7_6t_L U1144 ( .A(n818), .B(n817), .Y(n838) );
  XOR2xp5r_ASAP7_6t_L U1145 ( .A(n798), .B(n852), .Y(n817) );
  XOR2xp5r_ASAP7_6t_L U1146 ( .A(n853), .B(n797), .Y(n852) );
  XOR2xp5r_ASAP7_6t_L U1147 ( .A(n854), .B(n815), .Y(n797) );
  INVx1_ASAP7_6t_L U1148 ( .A(n813), .Y(n815) );
  XOR2xp5r_ASAP7_6t_L U1149 ( .A(n855), .B(n816), .Y(n813) );
  XOR2xp5r_ASAP7_6t_L U1150 ( .A(n810), .B(n809), .Y(n816) );
  NOR2xp5_ASAP7_6t_L U1151 ( .A(n96), .B(n170), .Y(n809) );
  XOR2xp5r_ASAP7_6t_L U1152 ( .A(n808), .B(n807), .Y(n810) );
  NOR2xp5_ASAP7_6t_L U1153 ( .A(n100), .B(n146), .Y(n807) );
  INVx1_ASAP7_6t_L U1154 ( .A(b[11]), .Y(n146) );
  NOR2xp5_ASAP7_6t_L U1155 ( .A(n98), .B(n126), .Y(n808) );
  INVx1_ASAP7_6t_L U1156 ( .A(b[12]), .Y(n126) );
  NOR2xp5_ASAP7_6t_L U1157 ( .A(n856), .B(n857), .Y(n855) );
  XOR2xp5r_ASAP7_6t_L U1158 ( .A(n858), .B(n814), .Y(n854) );
  XOR2xp5r_ASAP7_6t_L U1159 ( .A(n811), .B(n859), .Y(n814) );
  NAND2xp5R_ASAP7_6t_L U1160 ( .A(a[4]), .B(b[8]), .Y(n859) );
  NAND2xp5R_ASAP7_6t_L U1161 ( .A(a[3]), .B(b[9]), .Y(n811) );
  NOR2xp5_ASAP7_6t_L U1162 ( .A(n392), .B(n296), .Y(n858) );
  NOR2xp5_ASAP7_6t_L U1163 ( .A(n285), .B(n311), .Y(n853) );
  AOI21xp25_ASAP7_6t_L U1164 ( .A1(n860), .A2(n861), .B(n862), .Y(n798) );
  NOR3x1f_ASAP7_6t_L U1165 ( .A(n861), .B(n258), .C(n497), .Y(n862) );
  OAI22xp5_ASAP7_6t_L U1166 ( .A1(n863), .A2(n864), .B1(n865), .B2(n866), .Y(
        n818) );
  AOI21xp25_ASAP7_6t_L U1167 ( .A1(n867), .A2(n868), .B(n869), .Y(n851) );
  NOR3x1f_ASAP7_6t_L U1168 ( .A(n867), .B(n392), .C(n311), .Y(n869) );
  XOR2xp5r_ASAP7_6t_L U1169 ( .A(n832), .B(n833), .Y(n836) );
  OAI22xp5_ASAP7_6t_L U1170 ( .A1(n870), .A2(n871), .B1(n872), .B2(n873), .Y(
        n833) );
  XOR2xp5r_ASAP7_6t_L U1171 ( .A(n874), .B(n820), .Y(n832) );
  AOI21xp25_ASAP7_6t_L U1172 ( .A1(n875), .A2(n876), .B(n877), .Y(n820) );
  NOR3x1f_ASAP7_6t_L U1173 ( .A(n876), .B(n250), .C(n472), .Y(n877) );
  XOR2xp5r_ASAP7_6t_L U1174 ( .A(n878), .B(n821), .Y(n874) );
  XOR2xp5r_ASAP7_6t_L U1175 ( .A(n879), .B(n826), .Y(n821) );
  XOR2xp5r_ASAP7_6t_L U1176 ( .A(n880), .B(n825), .Y(n826) );
  NOR2xp5_ASAP7_6t_L U1177 ( .A(n361), .B(n280), .Y(n825) );
  NAND2xp5R_ASAP7_6t_L U1178 ( .A(a[8]), .B(b[4]), .Y(n880) );
  XOR2xp5r_ASAP7_6t_L U1179 ( .A(n881), .B(n823), .Y(n879) );
  NAND2xp5R_ASAP7_6t_L U1180 ( .A(b[2]), .B(a[10]), .Y(n823) );
  NAND2xp5R_ASAP7_6t_L U1181 ( .A(b[3]), .B(a[9]), .Y(n881) );
  NOR2xp5_ASAP7_6t_L U1182 ( .A(n160), .B(n99), .Y(n878) );
  AOI21xp25_ASAP7_6t_L U1183 ( .A1(n882), .A2(n883), .B(n884), .Y(n842) );
  NOR3x1f_ASAP7_6t_L U1184 ( .A(n882), .B(n185), .C(n99), .Y(n884) );
  NOR2xp5_ASAP7_6t_L U1185 ( .A(n114), .B(n97), .Y(n849) );
  INVx1_ASAP7_6t_L U1186 ( .A(a[12]), .Y(n114) );
  AOI22xp25_ASAP7_6t_L U1187 ( .A1(n885), .A2(n886), .B1(n887), .B2(n888), .Y(
        n839) );
  AO21x1_ASAP7_6t_L U1188 ( .A1(n79), .A2(n78), .B(n889), .Y(c[68]) );
  NOR3x1f_ASAP7_6t_L U1189 ( .A(n79), .B(n160), .C(n97), .Y(n889) );
  OAI22xp5_ASAP7_6t_L U1190 ( .A1(n890), .A2(n891), .B1(n892), .B2(n893), .Y(
        n78) );
  INVx1_ASAP7_6t_L U1191 ( .A(n894), .Y(n893) );
  INVx1_ASAP7_6t_L U1192 ( .A(n891), .Y(n892) );
  XOR2xp5r_ASAP7_6t_L U1193 ( .A(n844), .B(n895), .Y(n79) );
  XOR2xp5r_ASAP7_6t_L U1194 ( .A(n896), .B(n845), .Y(n895) );
  XOR2xp5r_ASAP7_6t_L U1195 ( .A(n847), .B(n897), .Y(n845) );
  XOR2xp5r_ASAP7_6t_L U1196 ( .A(n886), .B(n885), .Y(n897) );
  INVx1_ASAP7_6t_L U1197 ( .A(n887), .Y(n885) );
  XOR2xp5r_ASAP7_6t_L U1198 ( .A(n898), .B(n888), .Y(n887) );
  XOR2xp5r_ASAP7_6t_L U1199 ( .A(n867), .B(n868), .Y(n888) );
  OAI22xp5_ASAP7_6t_L U1200 ( .A1(n899), .A2(n900), .B1(n901), .B2(n902), .Y(
        n868) );
  XOR2xp5r_ASAP7_6t_L U1201 ( .A(n903), .B(n863), .Y(n867) );
  AOI21xp25_ASAP7_6t_L U1202 ( .A1(n904), .A2(n905), .B(n906), .Y(n863) );
  NOR3x1f_ASAP7_6t_L U1203 ( .A(n905), .B(n258), .C(n96), .Y(n906) );
  XOR2xp5r_ASAP7_6t_L U1204 ( .A(n865), .B(n907), .Y(n903) );
  NAND2xp5R_ASAP7_6t_L U1205 ( .A(b[6]), .B(a[5]), .Y(n907) );
  INVx1_ASAP7_6t_L U1206 ( .A(n864), .Y(n865) );
  XOR2xp5r_ASAP7_6t_L U1207 ( .A(n908), .B(n861), .Y(n864) );
  XOR2xp5r_ASAP7_6t_L U1208 ( .A(n860), .B(n909), .Y(n861) );
  NAND2xp5R_ASAP7_6t_L U1209 ( .A(a[2]), .B(b[9]), .Y(n909) );
  XOR2xp5r_ASAP7_6t_L U1210 ( .A(n856), .B(n857), .Y(n860) );
  NAND2xp5R_ASAP7_6t_L U1211 ( .A(a[0]), .B(b[11]), .Y(n857) );
  NAND2xp5R_ASAP7_6t_L U1212 ( .A(a[1]), .B(b[10]), .Y(n856) );
  XOR2xp5r_ASAP7_6t_L U1213 ( .A(n910), .B(n866), .Y(n908) );
  NAND2xp5R_ASAP7_6t_L U1214 ( .A(b[7]), .B(a[4]), .Y(n866) );
  NAND2xp5R_ASAP7_6t_L U1215 ( .A(a[3]), .B(b[8]), .Y(n910) );
  AOI21xp25_ASAP7_6t_L U1216 ( .A1(n911), .A2(n912), .B(n913), .Y(n898) );
  NOR3x1f_ASAP7_6t_L U1217 ( .A(n911), .B(n433), .C(n311), .Y(n913) );
  INVx1_ASAP7_6t_L U1218 ( .A(n914), .Y(n911) );
  XOR2xp5r_ASAP7_6t_L U1219 ( .A(n882), .B(n883), .Y(n886) );
  OAI22xp5_ASAP7_6t_L U1220 ( .A1(n915), .A2(n916), .B1(n917), .B2(n918), .Y(
        n883) );
  INVx1_ASAP7_6t_L U1221 ( .A(n917), .Y(n916) );
  XOR2xp5r_ASAP7_6t_L U1222 ( .A(n919), .B(n870), .Y(n882) );
  AOI21xp25_ASAP7_6t_L U1223 ( .A1(n920), .A2(n921), .B(n922), .Y(n870) );
  NOR3x1f_ASAP7_6t_L U1224 ( .A(n921), .B(n280), .C(n472), .Y(n922) );
  XOR2xp5r_ASAP7_6t_L U1225 ( .A(n923), .B(n871), .Y(n919) );
  INVx1_ASAP7_6t_L U1226 ( .A(n872), .Y(n871) );
  XOR2xp5r_ASAP7_6t_L U1227 ( .A(n876), .B(n924), .Y(n872) );
  XOR2xp5r_ASAP7_6t_L U1228 ( .A(n925), .B(n873), .Y(n924) );
  NAND2xp5R_ASAP7_6t_L U1229 ( .A(b[2]), .B(a[9]), .Y(n873) );
  NOR2xp5_ASAP7_6t_L U1230 ( .A(n250), .B(n472), .Y(n925) );
  XOR2xp5r_ASAP7_6t_L U1231 ( .A(n926), .B(n875), .Y(n876) );
  NOR2xp5_ASAP7_6t_L U1232 ( .A(n361), .B(n285), .Y(n875) );
  NAND2xp5R_ASAP7_6t_L U1233 ( .A(a[7]), .B(b[4]), .Y(n926) );
  NOR2xp5_ASAP7_6t_L U1234 ( .A(n185), .B(n99), .Y(n923) );
  NOR2xp5_ASAP7_6t_L U1235 ( .A(n927), .B(n928), .Y(n847) );
  NOR3x1f_ASAP7_6t_L U1236 ( .A(n929), .B(n930), .C(n931), .Y(n928) );
  NOR3x1f_ASAP7_6t_L U1237 ( .A(n932), .B(n212), .C(n99), .Y(n927) );
  INVx1_ASAP7_6t_L U1238 ( .A(n929), .Y(n932) );
  NOR2xp5_ASAP7_6t_L U1239 ( .A(n160), .B(n97), .Y(n896) );
  INVx1_ASAP7_6t_L U1240 ( .A(a[11]), .Y(n160) );
  OA22x1_ASAP7_6t_L U1241 ( .A1(n933), .A2(n934), .B1(n935), .B2(n936), .Y(
        n844) );
  INVx1_ASAP7_6t_L U1242 ( .A(n935), .Y(n933) );
  AO21x1_ASAP7_6t_L U1243 ( .A1(n81), .A2(n80), .B(n937), .Y(c[67]) );
  NOR3x1f_ASAP7_6t_L U1244 ( .A(n81), .B(n185), .C(n97), .Y(n937) );
  OAI22xp5_ASAP7_6t_L U1245 ( .A1(n938), .A2(n939), .B1(n940), .B2(n941), .Y(
        n80) );
  INVx1_ASAP7_6t_L U1246 ( .A(n942), .Y(n941) );
  INVx1_ASAP7_6t_L U1247 ( .A(n940), .Y(n939) );
  XOR2xp5r_ASAP7_6t_L U1248 ( .A(n890), .B(n943), .Y(n81) );
  XOR2xp5r_ASAP7_6t_L U1249 ( .A(n944), .B(n891), .Y(n943) );
  XOR2xp5r_ASAP7_6t_L U1250 ( .A(n934), .B(n945), .Y(n891) );
  XOR2xp5r_ASAP7_6t_L U1251 ( .A(n894), .B(n935), .Y(n945) );
  XOR2xp5r_ASAP7_6t_L U1252 ( .A(n946), .B(n936), .Y(n935) );
  XOR2xp5r_ASAP7_6t_L U1253 ( .A(n914), .B(n912), .Y(n936) );
  OAI22xp5_ASAP7_6t_L U1254 ( .A1(n947), .A2(n948), .B1(n949), .B2(n950), .Y(
        n912) );
  INVx1_ASAP7_6t_L U1255 ( .A(n948), .Y(n949) );
  XOR2xp5r_ASAP7_6t_L U1256 ( .A(n951), .B(n899), .Y(n914) );
  AOI21xp25_ASAP7_6t_L U1257 ( .A1(n952), .A2(n953), .B(n954), .Y(n899) );
  NOR3x1f_ASAP7_6t_L U1258 ( .A(n953), .B(n96), .C(n296), .Y(n954) );
  XOR2xp5r_ASAP7_6t_L U1259 ( .A(n955), .B(n901), .Y(n951) );
  INVx1_ASAP7_6t_L U1260 ( .A(n900), .Y(n901) );
  XOR2xp5r_ASAP7_6t_L U1261 ( .A(n956), .B(n905), .Y(n900) );
  XOR2xp5r_ASAP7_6t_L U1262 ( .A(n957), .B(n904), .Y(n905) );
  NOR2xp5_ASAP7_6t_L U1263 ( .A(n98), .B(n170), .Y(n904) );
  INVx1_ASAP7_6t_L U1264 ( .A(b[10]), .Y(n170) );
  NAND2xp5R_ASAP7_6t_L U1265 ( .A(b[9]), .B(a[1]), .Y(n957) );
  XOR2xp5r_ASAP7_6t_L U1266 ( .A(n958), .B(n902), .Y(n956) );
  NAND2xp5R_ASAP7_6t_L U1267 ( .A(b[7]), .B(a[3]), .Y(n902) );
  NAND2xp5R_ASAP7_6t_L U1268 ( .A(a[2]), .B(b[8]), .Y(n958) );
  NOR2xp5_ASAP7_6t_L U1269 ( .A(n433), .B(n311), .Y(n955) );
  AOI21xp25_ASAP7_6t_L U1270 ( .A1(n959), .A2(n960), .B(n961), .Y(n946) );
  NOR3x1f_ASAP7_6t_L U1271 ( .A(n959), .B(n433), .C(n361), .Y(n961) );
  NOR3x1f_ASAP7_6t_L U1272 ( .A(n962), .B(n212), .C(n97), .Y(n894) );
  XOR2xp5r_ASAP7_6t_L U1273 ( .A(n963), .B(n929), .Y(n934) );
  XOR2xp5r_ASAP7_6t_L U1274 ( .A(n964), .B(n915), .Y(n929) );
  AOI21xp25_ASAP7_6t_L U1275 ( .A1(n965), .A2(n966), .B(n967), .Y(n915) );
  NOR3x1f_ASAP7_6t_L U1276 ( .A(n966), .B(n280), .C(n537), .Y(n967) );
  XOR2xp5r_ASAP7_6t_L U1277 ( .A(n968), .B(n917), .Y(n964) );
  XOR2xp5r_ASAP7_6t_L U1278 ( .A(n921), .B(n969), .Y(n917) );
  XOR2xp5r_ASAP7_6t_L U1279 ( .A(n970), .B(n918), .Y(n969) );
  NAND2xp5R_ASAP7_6t_L U1280 ( .A(b[2]), .B(a[8]), .Y(n918) );
  NOR2xp5_ASAP7_6t_L U1281 ( .A(n280), .B(n472), .Y(n970) );
  XOR2xp5r_ASAP7_6t_L U1282 ( .A(n971), .B(n920), .Y(n921) );
  NOR2xp5_ASAP7_6t_L U1283 ( .A(n361), .B(n392), .Y(n920) );
  NAND2xp5R_ASAP7_6t_L U1284 ( .A(a[6]), .B(b[4]), .Y(n971) );
  NOR2xp5_ASAP7_6t_L U1285 ( .A(n212), .B(n99), .Y(n968) );
  INVx1_ASAP7_6t_L U1286 ( .A(a[9]), .Y(n212) );
  NOR2xp5_ASAP7_6t_L U1287 ( .A(n931), .B(n930), .Y(n963) );
  NOR2xp5_ASAP7_6t_L U1288 ( .A(n185), .B(n97), .Y(n944) );
  INVx1_ASAP7_6t_L U1289 ( .A(a[10]), .Y(n185) );
  AOI22xp25_ASAP7_6t_L U1290 ( .A1(n972), .A2(n962), .B1(n973), .B2(n974), .Y(
        n890) );
  NOR2xp5_ASAP7_6t_L U1291 ( .A(n83), .B(n82), .Y(c[66]) );
  XOR2xp5r_ASAP7_6t_L U1292 ( .A(n938), .B(n940), .Y(n82) );
  XOR2xp5r_ASAP7_6t_L U1293 ( .A(n962), .B(n975), .Y(n940) );
  XOR2xp5r_ASAP7_6t_L U1294 ( .A(n942), .B(n972), .Y(n975) );
  INVx1_ASAP7_6t_L U1295 ( .A(n973), .Y(n972) );
  XOR2xp5r_ASAP7_6t_L U1296 ( .A(n976), .B(n974), .Y(n973) );
  XOR2xp5r_ASAP7_6t_L U1297 ( .A(n959), .B(n960), .Y(n974) );
  AO22x1_ASAP7_6t_L U1298 ( .A1(n977), .A2(n978), .B1(n979), .B2(n980), .Y(
        n960) );
  INVx1_ASAP7_6t_L U1299 ( .A(n978), .Y(n979) );
  XOR2xp5r_ASAP7_6t_L U1300 ( .A(n981), .B(n947), .Y(n959) );
  AOI21xp25_ASAP7_6t_L U1301 ( .A1(n982), .A2(n983), .B(n984), .Y(n947) );
  NOR3x1f_ASAP7_6t_L U1302 ( .A(n983), .B(n96), .C(n311), .Y(n984) );
  XOR2xp5r_ASAP7_6t_L U1303 ( .A(n985), .B(n948), .Y(n981) );
  XOR2xp5r_ASAP7_6t_L U1304 ( .A(n986), .B(n953), .Y(n948) );
  XOR2xp5r_ASAP7_6t_L U1305 ( .A(n987), .B(n952), .Y(n953) );
  NOR2xp5_ASAP7_6t_L U1306 ( .A(n98), .B(n195), .Y(n952) );
  INVx1_ASAP7_6t_L U1307 ( .A(b[9]), .Y(n195) );
  NAND2xp5R_ASAP7_6t_L U1308 ( .A(b[8]), .B(a[1]), .Y(n987) );
  XOR2xp5r_ASAP7_6t_L U1309 ( .A(n988), .B(n950), .Y(n986) );
  NAND2xp5R_ASAP7_6t_L U1310 ( .A(b[6]), .B(a[3]), .Y(n950) );
  NAND2xp5R_ASAP7_6t_L U1311 ( .A(b[7]), .B(a[2]), .Y(n988) );
  NOR2xp5_ASAP7_6t_L U1312 ( .A(n433), .B(n361), .Y(n985) );
  AOI21xp25_ASAP7_6t_L U1313 ( .A1(n989), .A2(n990), .B(n991), .Y(n976) );
  NOR3x1f_ASAP7_6t_L U1314 ( .A(n989), .B(n433), .C(n417), .Y(n991) );
  NOR3x1f_ASAP7_6t_L U1315 ( .A(n992), .B(n285), .C(n537), .Y(n942) );
  INVx1_ASAP7_6t_L U1316 ( .A(a[6]), .Y(n285) );
  INVx1_ASAP7_6t_L U1317 ( .A(n993), .Y(n962) );
  XOR2xp5r_ASAP7_6t_L U1318 ( .A(n930), .B(n994), .Y(n993) );
  NAND2xp5R_ASAP7_6t_L U1319 ( .A(b[0]), .B(a[9]), .Y(n994) );
  XOR2xp5r_ASAP7_6t_L U1320 ( .A(n966), .B(n995), .Y(n930) );
  XOR2xp5r_ASAP7_6t_L U1321 ( .A(n996), .B(n931), .Y(n995) );
  NAND2xp5R_ASAP7_6t_L U1322 ( .A(b[1]), .B(a[8]), .Y(n931) );
  NOR2xp5_ASAP7_6t_L U1323 ( .A(n280), .B(n537), .Y(n996) );
  XOR2xp5r_ASAP7_6t_L U1324 ( .A(n997), .B(n965), .Y(n966) );
  NOR2xp5_ASAP7_6t_L U1325 ( .A(n417), .B(n392), .Y(n965) );
  NAND2xp5R_ASAP7_6t_L U1326 ( .A(a[6]), .B(b[3]), .Y(n997) );
  AOI22xp25_ASAP7_6t_L U1327 ( .A1(n998), .A2(n999), .B1(n1000), .B2(n1001), 
        .Y(n938) );
  AOI21xp25_ASAP7_6t_L U1328 ( .A1(n1002), .A2(n1003), .B(n1004), .Y(n83) );
  NOR3x1f_ASAP7_6t_L U1329 ( .A(n1002), .B(n280), .C(n99), .Y(n1004) );
  AO21x1_ASAP7_6t_L U1330 ( .A1(n85), .A2(n84), .B(n1005), .Y(c[65]) );
  NOR3x1f_ASAP7_6t_L U1331 ( .A(n85), .B(n250), .C(n97), .Y(n1005) );
  OAI22xp5_ASAP7_6t_L U1332 ( .A1(n1006), .A2(n1007), .B1(n1008), .B2(n1009), 
        .Y(n84) );
  XOR2xp5r_ASAP7_6t_L U1333 ( .A(n1003), .B(n1010), .Y(n85) );
  XOR2xp5r_ASAP7_6t_L U1334 ( .A(n1011), .B(n1002), .Y(n1010) );
  XOR2xp5r_ASAP7_6t_L U1335 ( .A(n999), .B(n1012), .Y(n1002) );
  XOR2xp5r_ASAP7_6t_L U1336 ( .A(n1013), .B(n998), .Y(n1012) );
  INVx1_ASAP7_6t_L U1337 ( .A(n1000), .Y(n998) );
  XOR2xp5r_ASAP7_6t_L U1338 ( .A(n1014), .B(n1001), .Y(n1000) );
  XOR2xp5r_ASAP7_6t_L U1339 ( .A(n990), .B(n989), .Y(n1001) );
  XOR2xp5r_ASAP7_6t_L U1340 ( .A(n1015), .B(n977), .Y(n989) );
  AO21x1_ASAP7_6t_L U1341 ( .A1(n1016), .A2(n1017), .B(n1018), .Y(n977) );
  NOR3x1f_ASAP7_6t_L U1342 ( .A(n1017), .B(n96), .C(n361), .Y(n1018) );
  XOR2xp5r_ASAP7_6t_L U1343 ( .A(n1019), .B(n978), .Y(n1015) );
  XOR2xp5r_ASAP7_6t_L U1344 ( .A(n983), .B(n1020), .Y(n978) );
  XOR2xp5r_ASAP7_6t_L U1345 ( .A(n980), .B(n1021), .Y(n1020) );
  NAND2xp5R_ASAP7_6t_L U1346 ( .A(b[6]), .B(a[2]), .Y(n1021) );
  NOR2xp5_ASAP7_6t_L U1347 ( .A(n361), .B(n497), .Y(n980) );
  INVx1_ASAP7_6t_L U1348 ( .A(b[5]), .Y(n361) );
  XOR2xp5r_ASAP7_6t_L U1349 ( .A(n1022), .B(n982), .Y(n983) );
  NOR2xp5_ASAP7_6t_L U1350 ( .A(n98), .B(n258), .Y(n982) );
  INVx1_ASAP7_6t_L U1351 ( .A(b[8]), .Y(n258) );
  NAND2xp5R_ASAP7_6t_L U1352 ( .A(a[1]), .B(b[7]), .Y(n1022) );
  NOR2xp5_ASAP7_6t_L U1353 ( .A(n433), .B(n417), .Y(n1019) );
  OAI22xp5_ASAP7_6t_L U1354 ( .A1(n1023), .A2(n1024), .B1(n1025), .B2(n1026), 
        .Y(n990) );
  NOR2xp5_ASAP7_6t_L U1355 ( .A(n1027), .B(n1028), .Y(n1014) );
  NOR3x1f_ASAP7_6t_L U1356 ( .A(n1029), .B(n1030), .C(n1031), .Y(n1028) );
  NOR3x1f_ASAP7_6t_L U1357 ( .A(n1032), .B(n433), .C(n472), .Y(n1027) );
  NOR2xp5_ASAP7_6t_L U1358 ( .A(n280), .B(n99), .Y(n1013) );
  XOR2xp5r_ASAP7_6t_L U1359 ( .A(n1033), .B(n992), .Y(n999) );
  NAND2xp5R_ASAP7_6t_L U1360 ( .A(b[3]), .B(a[5]), .Y(n992) );
  NAND2xp5R_ASAP7_6t_L U1361 ( .A(a[6]), .B(b[2]), .Y(n1033) );
  NOR2xp5_ASAP7_6t_L U1362 ( .A(n250), .B(n97), .Y(n1011) );
  INVx1_ASAP7_6t_L U1363 ( .A(a[8]), .Y(n250) );
  AO21x1_ASAP7_6t_L U1364 ( .A1(n1034), .A2(n1035), .B(n1036), .Y(n1003) );
  NOR3x1f_ASAP7_6t_L U1365 ( .A(n1035), .B(n392), .C(n537), .Y(n1036) );
  AO21x1_ASAP7_6t_L U1366 ( .A1(n87), .A2(n86), .B(n1037), .Y(c[64]) );
  NOR3x1f_ASAP7_6t_L U1367 ( .A(n87), .B(n280), .C(n97), .Y(n1037) );
  OAI22xp5_ASAP7_6t_L U1368 ( .A1(n1038), .A2(n1039), .B1(n1040), .B2(n1041), 
        .Y(n86) );
  INVx1_ASAP7_6t_L U1369 ( .A(n1040), .Y(n1039) );
  XOR2xp5r_ASAP7_6t_L U1370 ( .A(n1042), .B(n1043), .Y(n87) );
  XOR2xp5r_ASAP7_6t_L U1371 ( .A(n1044), .B(n1008), .Y(n1043) );
  INVx1_ASAP7_6t_L U1372 ( .A(n1007), .Y(n1008) );
  XOR2xp5r_ASAP7_6t_L U1373 ( .A(n1045), .B(n1035), .Y(n1007) );
  XOR2xp5r_ASAP7_6t_L U1374 ( .A(n1046), .B(n1034), .Y(n1035) );
  XOR2xp5r_ASAP7_6t_L U1375 ( .A(n1047), .B(n1032), .Y(n1034) );
  INVx1_ASAP7_6t_L U1376 ( .A(n1029), .Y(n1032) );
  XOR2xp5r_ASAP7_6t_L U1377 ( .A(n1048), .B(n1023), .Y(n1029) );
  AOI21xp25_ASAP7_6t_L U1378 ( .A1(n1049), .A2(n1050), .B(n1051), .Y(n1023) );
  NOR3x1f_ASAP7_6t_L U1379 ( .A(n1050), .B(n96), .C(n417), .Y(n1051) );
  XOR2xp5r_ASAP7_6t_L U1380 ( .A(n1052), .B(n1025), .Y(n1048) );
  INVx1_ASAP7_6t_L U1381 ( .A(n1024), .Y(n1025) );
  XOR2xp5r_ASAP7_6t_L U1382 ( .A(n1017), .B(n1053), .Y(n1024) );
  XOR2xp5r_ASAP7_6t_L U1383 ( .A(n1026), .B(n1054), .Y(n1053) );
  NAND2xp5R_ASAP7_6t_L U1384 ( .A(b[5]), .B(a[2]), .Y(n1054) );
  NAND2xp5R_ASAP7_6t_L U1385 ( .A(b[4]), .B(a[3]), .Y(n1026) );
  XOR2xp5r_ASAP7_6t_L U1386 ( .A(n1055), .B(n1016), .Y(n1017) );
  NOR2xp5_ASAP7_6t_L U1387 ( .A(n98), .B(n296), .Y(n1016) );
  INVx1_ASAP7_6t_L U1388 ( .A(b[7]), .Y(n296) );
  NAND2xp5R_ASAP7_6t_L U1389 ( .A(a[1]), .B(b[6]), .Y(n1055) );
  NOR2xp5_ASAP7_6t_L U1390 ( .A(n433), .B(n472), .Y(n1052) );
  NOR2xp5_ASAP7_6t_L U1391 ( .A(n1031), .B(n1030), .Y(n1047) );
  INVx1_ASAP7_6t_L U1392 ( .A(n1056), .Y(n1030) );
  OR2x2_ASAP7_6t_L U1393 ( .A(n1057), .B(n1058), .Y(n1046) );
  XOR2xp5r_ASAP7_6t_L U1394 ( .A(n1059), .B(n1009), .Y(n1045) );
  NAND2xp5R_ASAP7_6t_L U1395 ( .A(b[1]), .B(a[6]), .Y(n1009) );
  NAND2xp5R_ASAP7_6t_L U1396 ( .A(b[2]), .B(a[5]), .Y(n1059) );
  NOR2xp5_ASAP7_6t_L U1397 ( .A(n280), .B(n97), .Y(n1044) );
  INVx1_ASAP7_6t_L U1398 ( .A(a[7]), .Y(n280) );
  INVx1_ASAP7_6t_L U1399 ( .A(n1006), .Y(n1042) );
  AOI21xp25_ASAP7_6t_L U1400 ( .A1(n1058), .A2(n1060), .B(n1061), .Y(n1006) );
  NOR3x1f_ASAP7_6t_L U1401 ( .A(n1060), .B(n392), .C(n99), .Y(n1061) );
  NOR2xp5_ASAP7_6t_L U1402 ( .A(n88), .B(n89), .Y(c[63]) );
  XOR2xp5r_ASAP7_6t_L U1403 ( .A(n1038), .B(n1040), .Y(n89) );
  XOR2xp5r_ASAP7_6t_L U1404 ( .A(n1060), .B(n1062), .Y(n1040) );
  XOR2xp5r_ASAP7_6t_L U1405 ( .A(n1063), .B(n1041), .Y(n1062) );
  NAND2xp5R_ASAP7_6t_L U1406 ( .A(b[0]), .B(a[6]), .Y(n1041) );
  NOR2xp5_ASAP7_6t_L U1407 ( .A(n392), .B(n99), .Y(n1063) );
  XOR2xp5r_ASAP7_6t_L U1408 ( .A(n1064), .B(n1058), .Y(n1060) );
  XOR2xp5r_ASAP7_6t_L U1409 ( .A(n1056), .B(n1057), .Y(n1058) );
  NAND2xp5R_ASAP7_6t_L U1410 ( .A(b[2]), .B(a[4]), .Y(n1057) );
  XOR2xp5r_ASAP7_6t_L U1411 ( .A(n1065), .B(n1050), .Y(n1056) );
  XOR2xp5r_ASAP7_6t_L U1412 ( .A(n1066), .B(n1049), .Y(n1050) );
  NOR2xp5_ASAP7_6t_L U1413 ( .A(n311), .B(n98), .Y(n1049) );
  INVx1_ASAP7_6t_L U1414 ( .A(b[6]), .Y(n311) );
  NAND2xp5R_ASAP7_6t_L U1415 ( .A(a[1]), .B(b[5]), .Y(n1066) );
  XOR2xp5r_ASAP7_6t_L U1416 ( .A(n1067), .B(n1031), .Y(n1065) );
  NAND2xp5R_ASAP7_6t_L U1417 ( .A(b[3]), .B(a[3]), .Y(n1031) );
  NAND2xp5R_ASAP7_6t_L U1418 ( .A(b[4]), .B(a[2]), .Y(n1067) );
  OR2x2_ASAP7_6t_L U1419 ( .A(n1068), .B(n1069), .Y(n1064) );
  AOI21xp25_ASAP7_6t_L U1420 ( .A1(n1070), .A2(n1071), .B(n1072), .Y(n1038) );
  NOR3x1f_ASAP7_6t_L U1421 ( .A(n1071), .B(n497), .C(n537), .Y(n1072) );
  INVx1_ASAP7_6t_L U1422 ( .A(a[3]), .Y(n497) );
  AOI22xp25_ASAP7_6t_L U1423 ( .A1(n1073), .A2(n1074), .B1(n1075), .B2(n1076), 
        .Y(n88) );
  AO21x1_ASAP7_6t_L U1424 ( .A1(n90), .A2(n91), .B(n1077), .Y(c[62]) );
  NOR3x1f_ASAP7_6t_L U1425 ( .A(n90), .B(n392), .C(n97), .Y(n1077) );
  INVx1_ASAP7_6t_L U1426 ( .A(a[5]), .Y(n392) );
  OAI22xp5_ASAP7_6t_L U1427 ( .A1(n1078), .A2(n1079), .B1(n1080), .B2(n1081), 
        .Y(n91) );
  INVx1_ASAP7_6t_L U1428 ( .A(n1079), .Y(n1080) );
  XOR2xp5r_ASAP7_6t_L U1429 ( .A(n1082), .B(n1073), .Y(n90) );
  AO21x1_ASAP7_6t_L U1430 ( .A1(n1083), .A2(n1084), .B(n1085), .Y(n1073) );
  NOR3x1f_ASAP7_6t_L U1431 ( .A(n1084), .B(n96), .C(n537), .Y(n1085) );
  INVx1_ASAP7_6t_L U1432 ( .A(b[2]), .Y(n537) );
  XOR2xp5r_ASAP7_6t_L U1433 ( .A(n1075), .B(n1086), .Y(n1082) );
  NAND2xp5R_ASAP7_6t_L U1434 ( .A(b[0]), .B(a[5]), .Y(n1086) );
  INVx1_ASAP7_6t_L U1435 ( .A(n1074), .Y(n1075) );
  XOR2xp5r_ASAP7_6t_L U1436 ( .A(n1087), .B(n1071), .Y(n1074) );
  XOR2xp5r_ASAP7_6t_L U1437 ( .A(n1070), .B(n1088), .Y(n1071) );
  NAND2xp5R_ASAP7_6t_L U1438 ( .A(b[3]), .B(a[2]), .Y(n1088) );
  XOR2xp5r_ASAP7_6t_L U1439 ( .A(n1069), .B(n1068), .Y(n1070) );
  NAND2xp5R_ASAP7_6t_L U1440 ( .A(b[4]), .B(a[1]), .Y(n1068) );
  NAND2xp5R_ASAP7_6t_L U1441 ( .A(b[5]), .B(a[0]), .Y(n1069) );
  XOR2xp5r_ASAP7_6t_L U1442 ( .A(n1089), .B(n1076), .Y(n1087) );
  NOR2xp5_ASAP7_6t_L U1443 ( .A(n99), .B(n433), .Y(n1076) );
  NAND2xp5R_ASAP7_6t_L U1444 ( .A(b[2]), .B(a[3]), .Y(n1089) );
  AO21x1_ASAP7_6t_L U1445 ( .A1(n92), .A2(n93), .B(n1090), .Y(c[61]) );
  NOR3x1f_ASAP7_6t_L U1446 ( .A(n93), .B(n433), .C(n97), .Y(n1090) );
  XOR2xp5r_ASAP7_6t_L U1447 ( .A(n1091), .B(n1078), .Y(n93) );
  AOI21xp25_ASAP7_6t_L U1448 ( .A1(n1092), .A2(n1093), .B(n1094), .Y(n1078) );
  NOR3x1f_ASAP7_6t_L U1449 ( .A(n1093), .B(n96), .C(n99), .Y(n1094) );
  XOR2xp5r_ASAP7_6t_L U1450 ( .A(n1095), .B(n1079), .Y(n1091) );
  XOR2xp5r_ASAP7_6t_L U1451 ( .A(n1096), .B(n1084), .Y(n1079) );
  XOR2xp5r_ASAP7_6t_L U1452 ( .A(n1083), .B(n1097), .Y(n1084) );
  NAND2xp5R_ASAP7_6t_L U1453 ( .A(b[3]), .B(a[1]), .Y(n1097) );
  NOR2xp5_ASAP7_6t_L U1454 ( .A(n417), .B(n98), .Y(n1083) );
  INVx1_ASAP7_6t_L U1455 ( .A(b[4]), .Y(n417) );
  XOR2xp5r_ASAP7_6t_L U1456 ( .A(n1098), .B(n1081), .Y(n1096) );
  NAND2xp5R_ASAP7_6t_L U1457 ( .A(b[1]), .B(a[3]), .Y(n1081) );
  NAND2xp5R_ASAP7_6t_L U1458 ( .A(b[2]), .B(a[2]), .Y(n1098) );
  NOR2xp5_ASAP7_6t_L U1459 ( .A(n433), .B(n97), .Y(n1095) );
  INVx1_ASAP7_6t_L U1460 ( .A(b[0]), .Y(n97) );
  INVx1_ASAP7_6t_L U1461 ( .A(a[4]), .Y(n433) );
  NOR2xp5_ASAP7_6t_L U1462 ( .A(n1099), .B(n1158), .Y(n92) );
  XOR2xp5r_ASAP7_6t_L U1463 ( .A(n1100), .B(n1093), .Y(n1158) );
  XOR2xp5r_ASAP7_6t_L U1464 ( .A(n1101), .B(n1092), .Y(n1093) );
  NOR2xp5_ASAP7_6t_L U1465 ( .A(n472), .B(n98), .Y(n1092) );
  INVx1_ASAP7_6t_L U1466 ( .A(a[0]), .Y(n98) );
  INVx1_ASAP7_6t_L U1467 ( .A(b[3]), .Y(n472) );
  NAND2xp5R_ASAP7_6t_L U1468 ( .A(a[1]), .B(b[2]), .Y(n1101) );
  XOR2xp5r_ASAP7_6t_L U1469 ( .A(n1102), .B(n1099), .Y(n1100) );
  NOR2xp5_ASAP7_6t_L U1470 ( .A(n99), .B(n96), .Y(n1102) );
  INVx1_ASAP7_6t_L U1471 ( .A(a[2]), .Y(n96) );
  NAND2xp5R_ASAP7_6t_L U1472 ( .A(b[0]), .B(a[3]), .Y(n1099) );
  NOR3x1f_ASAP7_6t_L U1473 ( .A(n95), .B(n100), .C(n99), .Y(c[59]) );
  INVx1_ASAP7_6t_L U1474 ( .A(b[1]), .Y(n99) );
  INVx1_ASAP7_6t_L U1475 ( .A(a[1]), .Y(n100) );
  NAND2xp5R_ASAP7_6t_L U1476 ( .A(b[2]), .B(a[0]), .Y(n95) );
endmodule

