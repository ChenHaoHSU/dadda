
module DADDA_16x16 ( a, b, out );
  input [15:0] a;
  input [15:0] b;
  output [31:0] out;
  wire   c_182_, add_290_CI, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1007, n1009, n1011, n1013, n1015, n1017, n1019, n1021,
         n1023, n1025, n1027, n1029, n1031, n1033, n1035, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1054, n1055, n1057, n1058, n1060, n1061, n1063,
         n1064, n1066, n1067, n1069, n1070, n1072, n1073, n1075, n1076, n1078,
         n1079, n1081, n1082, n1084, n1085, n1087, n1088, n1090, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151;
  wire   [255:1] p;
  wire   [209:182] s;

  FAxp33_ASAP7_6t_L add_290_U1_0 ( .A(p[1]), .B(p[16]), .CI(add_290_CI), .CON(
        n1093), .SN(n1092) );
  FAxp33_ASAP7_6t_L add_290_U1_1 ( .A(s[182]), .B(p[32]), .CI(n1090), .CON(
        n1095), .SN(n1094) );
  FAxp33_ASAP7_6t_L add_290_U1_2 ( .A(c_182_), .B(s[183]), .CI(n1088), .CON(
        n1097), .SN(n1096) );
  FAxp33_ASAP7_6t_L add_290_U1_3 ( .A(n1087), .B(s[184]), .CI(n1085), .CON(
        n1099), .SN(n1098) );
  FAxp33_ASAP7_6t_L add_290_U1_4 ( .A(n1084), .B(s[185]), .CI(n1082), .CON(
        n1101), .SN(n1100) );
  FAxp33_ASAP7_6t_L add_290_U1_5 ( .A(n1081), .B(s[186]), .CI(n1079), .CON(
        n1103), .SN(n1102) );
  FAxp33_ASAP7_6t_L add_290_U1_6 ( .A(n1078), .B(s[187]), .CI(n1076), .CON(
        n1105), .SN(n1104) );
  FAxp33_ASAP7_6t_L add_290_U1_7 ( .A(n1075), .B(s[188]), .CI(n1073), .CON(
        n1107), .SN(n1106) );
  FAxp33_ASAP7_6t_L add_290_U1_8 ( .A(n1072), .B(s[189]), .CI(n1070), .CON(
        n1109), .SN(n1108) );
  FAxp33_ASAP7_6t_L add_290_U1_9 ( .A(n1069), .B(s[190]), .CI(n1067), .CON(
        n1111), .SN(n1110) );
  FAxp33_ASAP7_6t_L add_290_U1_10 ( .A(n1066), .B(s[191]), .CI(n1064), .CON(
        n1113), .SN(n1112) );
  FAxp33_ASAP7_6t_L add_290_U1_11 ( .A(n1063), .B(s[192]), .CI(n1061), .CON(
        n1115), .SN(n1114) );
  FAxp33_ASAP7_6t_L add_290_U1_12 ( .A(n1060), .B(s[193]), .CI(n1058), .CON(
        n1117), .SN(n1116) );
  FAxp33_ASAP7_6t_L add_290_U1_13 ( .A(n1057), .B(s[194]), .CI(n1055), .CON(
        n1119), .SN(n1118) );
  FAxp33_ASAP7_6t_L add_290_U1_14 ( .A(n1054), .B(s[195]), .CI(n1052), .CON(
        n1121), .SN(n1120) );
  FAxp33_ASAP7_6t_L add_290_U1_15 ( .A(n1037), .B(s[196]), .CI(n1035), .CON(
        n1123), .SN(n1122) );
  FAxp33_ASAP7_6t_L add_290_U1_16 ( .A(n1039), .B(s[197]), .CI(n1033), .CON(
        n1125), .SN(n1124) );
  FAxp33_ASAP7_6t_L add_290_U1_17 ( .A(n1038), .B(s[198]), .CI(n1031), .CON(
        n1127), .SN(n1126) );
  FAxp33_ASAP7_6t_L add_290_U1_18 ( .A(n1040), .B(s[199]), .CI(n1029), .CON(
        n1129), .SN(n1128) );
  FAxp33_ASAP7_6t_L add_290_U1_19 ( .A(n1041), .B(s[200]), .CI(n1027), .CON(
        n1131), .SN(n1130) );
  FAxp33_ASAP7_6t_L add_290_U1_20 ( .A(n1042), .B(s[201]), .CI(n1025), .CON(
        n1133), .SN(n1132) );
  FAxp33_ASAP7_6t_L add_290_U1_21 ( .A(n1043), .B(s[202]), .CI(n1023), .CON(
        n1135), .SN(n1134) );
  FAxp33_ASAP7_6t_L add_290_U1_22 ( .A(n1044), .B(s[203]), .CI(n1021), .CON(
        n1137), .SN(n1136) );
  FAxp33_ASAP7_6t_L add_290_U1_23 ( .A(n1045), .B(s[204]), .CI(n1019), .CON(
        n1139), .SN(n1138) );
  FAxp33_ASAP7_6t_L add_290_U1_24 ( .A(n1046), .B(s[205]), .CI(n1017), .CON(
        n1141), .SN(n1140) );
  FAxp33_ASAP7_6t_L add_290_U1_25 ( .A(n1047), .B(s[206]), .CI(n1015), .CON(
        n1143), .SN(n1142) );
  FAxp33_ASAP7_6t_L add_290_U1_26 ( .A(n1048), .B(s[207]), .CI(n1013), .CON(
        n1145), .SN(n1144) );
  FAxp33_ASAP7_6t_L add_290_U1_27 ( .A(n1049), .B(s[208]), .CI(n1011), .CON(
        n1147), .SN(n1146) );
  FAxp33_ASAP7_6t_L add_290_U1_28 ( .A(n1050), .B(s[209]), .CI(n1009), .CON(
        n1149), .SN(n1148) );
  FAxp33_ASAP7_6t_L add_290_U1_29 ( .A(n1051), .B(p[255]), .CI(n1007), .CON(
        n1151), .SN(n1150) );
  TIELOxp5_ASAP7_6t_L U291 ( .L(add_290_CI) );
  XOR2xp5r_ASAP7_6t_L U292 ( .A(n35), .B(n36), .Y(s[209]) );
  NAND2xp5R_ASAP7_6t_L U293 ( .A(a[15]), .B(b[14]), .Y(n35) );
  XOR2xp5r_ASAP7_6t_L U294 ( .A(n37), .B(n38), .Y(s[208]) );
  NAND2xp5R_ASAP7_6t_L U295 ( .A(a[15]), .B(b[13]), .Y(n37) );
  XOR2xp5r_ASAP7_6t_L U296 ( .A(n39), .B(n40), .Y(s[207]) );
  NOR2xp5_ASAP7_6t_L U297 ( .A(n41), .B(n42), .Y(n39) );
  XOR2xp5r_ASAP7_6t_L U298 ( .A(n43), .B(n44), .Y(s[206]) );
  XOR2xp5r_ASAP7_6t_L U299 ( .A(n45), .B(n46), .Y(s[205]) );
  XOR2xp5r_ASAP7_6t_L U300 ( .A(n47), .B(n48), .Y(s[204]) );
  XOR2xp5r_ASAP7_6t_L U301 ( .A(n49), .B(n50), .Y(s[203]) );
  XOR2xp5r_ASAP7_6t_L U302 ( .A(n51), .B(n52), .Y(s[202]) );
  XOR2xp5r_ASAP7_6t_L U303 ( .A(n53), .B(n54), .Y(s[201]) );
  XOR2xp5r_ASAP7_6t_L U304 ( .A(n55), .B(n56), .Y(s[200]) );
  XOR2xp5r_ASAP7_6t_L U305 ( .A(n57), .B(n58), .Y(s[199]) );
  XOR2xp5r_ASAP7_6t_L U306 ( .A(n59), .B(n60), .Y(s[198]) );
  XOR2xp5r_ASAP7_6t_L U307 ( .A(n61), .B(n62), .Y(s[197]) );
  XOR2xp5r_ASAP7_6t_L U308 ( .A(n63), .B(n64), .Y(s[196]) );
  XOR2xp5r_ASAP7_6t_L U309 ( .A(n65), .B(n66), .Y(s[195]) );
  XOR2xp5r_ASAP7_6t_L U310 ( .A(n67), .B(n68), .Y(s[194]) );
  XOR2xp5r_ASAP7_6t_L U311 ( .A(n69), .B(n70), .Y(s[193]) );
  XOR2xp5r_ASAP7_6t_L U312 ( .A(n71), .B(n72), .Y(s[192]) );
  XOR2xp5r_ASAP7_6t_L U313 ( .A(n73), .B(n74), .Y(s[191]) );
  XOR2xp5r_ASAP7_6t_L U314 ( .A(n75), .B(n76), .Y(s[190]) );
  XOR2xp5r_ASAP7_6t_L U315 ( .A(n77), .B(n78), .Y(s[189]) );
  XOR2xp5r_ASAP7_6t_L U316 ( .A(n79), .B(n80), .Y(s[188]) );
  XOR2xp5r_ASAP7_6t_L U317 ( .A(n81), .B(n82), .Y(s[187]) );
  XOR2xp5r_ASAP7_6t_L U318 ( .A(n83), .B(n84), .Y(s[186]) );
  XOR2xp5r_ASAP7_6t_L U319 ( .A(n85), .B(n86), .Y(s[185]) );
  NAND2xp5R_ASAP7_6t_L U320 ( .A(a[5]), .B(b[0]), .Y(n85) );
  XOR2xp5r_ASAP7_6t_L U321 ( .A(n87), .B(n88), .Y(s[184]) );
  NOR2xp5_ASAP7_6t_L U322 ( .A(n89), .B(n90), .Y(n87) );
  XOR2xp5r_ASAP7_6t_L U323 ( .A(n91), .B(n92), .Y(s[183]) );
  NAND2xp5R_ASAP7_6t_L U324 ( .A(b[0]), .B(a[3]), .Y(n92) );
  XOR2xp5r_ASAP7_6t_L U325 ( .A(n93), .B(n94), .Y(s[182]) );
  NAND2xp5R_ASAP7_6t_L U326 ( .A(b[1]), .B(a[1]), .Y(n93) );
  NOR2xp5_ASAP7_6t_L U327 ( .A(n95), .B(n90), .Y(p[32]) );
  NOR2xp5_ASAP7_6t_L U328 ( .A(n41), .B(n96), .Y(p[255]) );
  NOR2xp5_ASAP7_6t_L U329 ( .A(n97), .B(n98), .Y(p[1]) );
  NOR2xp5_ASAP7_6t_L U330 ( .A(n99), .B(n90), .Y(p[16]) );
  NOR2xp5_ASAP7_6t_L U331 ( .A(n97), .B(n90), .Y(out[0]) );
  INVx1_ASAP7_6t_L U332 ( .A(n1151), .Y(out[31]) );
  INVx1_ASAP7_6t_L U333 ( .A(n1150), .Y(out[30]) );
  INVx1_ASAP7_6t_L U334 ( .A(n1149), .Y(n1007) );
  INVx1_ASAP7_6t_L U335 ( .A(n1148), .Y(out[29]) );
  INVx1_ASAP7_6t_L U336 ( .A(n1147), .Y(n1009) );
  INVx1_ASAP7_6t_L U337 ( .A(n1146), .Y(out[28]) );
  INVx1_ASAP7_6t_L U338 ( .A(n1145), .Y(n1011) );
  INVx1_ASAP7_6t_L U339 ( .A(n1144), .Y(out[27]) );
  INVx1_ASAP7_6t_L U340 ( .A(n1143), .Y(n1013) );
  INVx1_ASAP7_6t_L U341 ( .A(n1142), .Y(out[26]) );
  INVx1_ASAP7_6t_L U342 ( .A(n1141), .Y(n1015) );
  INVx1_ASAP7_6t_L U343 ( .A(n1140), .Y(out[25]) );
  INVx1_ASAP7_6t_L U344 ( .A(n1139), .Y(n1017) );
  INVx1_ASAP7_6t_L U345 ( .A(n1138), .Y(out[24]) );
  INVx1_ASAP7_6t_L U346 ( .A(n1137), .Y(n1019) );
  INVx1_ASAP7_6t_L U347 ( .A(n1136), .Y(out[23]) );
  INVx1_ASAP7_6t_L U348 ( .A(n1135), .Y(n1021) );
  INVx1_ASAP7_6t_L U349 ( .A(n1134), .Y(out[22]) );
  INVx1_ASAP7_6t_L U350 ( .A(n1133), .Y(n1023) );
  INVx1_ASAP7_6t_L U351 ( .A(n1132), .Y(out[21]) );
  INVx1_ASAP7_6t_L U352 ( .A(n1131), .Y(n1025) );
  INVx1_ASAP7_6t_L U353 ( .A(n1130), .Y(out[20]) );
  INVx1_ASAP7_6t_L U354 ( .A(n1129), .Y(n1027) );
  INVx1_ASAP7_6t_L U355 ( .A(n1128), .Y(out[19]) );
  INVx1_ASAP7_6t_L U356 ( .A(n1127), .Y(n1029) );
  INVx1_ASAP7_6t_L U357 ( .A(n1126), .Y(out[18]) );
  INVx1_ASAP7_6t_L U358 ( .A(n1125), .Y(n1031) );
  INVx1_ASAP7_6t_L U359 ( .A(n1124), .Y(out[17]) );
  INVx1_ASAP7_6t_L U360 ( .A(n1123), .Y(n1033) );
  INVx1_ASAP7_6t_L U361 ( .A(n1122), .Y(out[16]) );
  INVx1_ASAP7_6t_L U362 ( .A(n1121), .Y(n1035) );
  INVx1_ASAP7_6t_L U363 ( .A(n1120), .Y(out[15]) );
  OAI22xp5_ASAP7_6t_L U364 ( .A1(n100), .A2(n101), .B1(n66), .B2(n65), .Y(
        n1037) );
  INVx1_ASAP7_6t_L U365 ( .A(n102), .Y(n65) );
  XOR2xp5r_ASAP7_6t_L U366 ( .A(n103), .B(n104), .Y(n102) );
  XOR2xp5r_ASAP7_6t_L U367 ( .A(n100), .B(n105), .Y(n66) );
  INVx1_ASAP7_6t_L U368 ( .A(n105), .Y(n101) );
  XOR2xp5r_ASAP7_6t_L U369 ( .A(n106), .B(n107), .Y(n105) );
  AOI22xp25_ASAP7_6t_L U370 ( .A1(n108), .A2(n109), .B1(n110), .B2(n111), .Y(
        n100) );
  OAI22xp5_ASAP7_6t_L U371 ( .A1(n112), .A2(n113), .B1(n61), .B2(n62), .Y(
        n1038) );
  XOR2xp5r_ASAP7_6t_L U372 ( .A(n114), .B(n112), .Y(n62) );
  XOR2xp5r_ASAP7_6t_L U373 ( .A(n115), .B(n116), .Y(n61) );
  INVx1_ASAP7_6t_L U374 ( .A(n117), .Y(n115) );
  INVx1_ASAP7_6t_L U375 ( .A(n114), .Y(n113) );
  XOR2xp5r_ASAP7_6t_L U376 ( .A(n118), .B(n119), .Y(n114) );
  AOI22xp25_ASAP7_6t_L U377 ( .A1(n120), .A2(n121), .B1(n122), .B2(n123), .Y(
        n112) );
  OAI22xp5_ASAP7_6t_L U378 ( .A1(n124), .A2(n125), .B1(n63), .B2(n64), .Y(
        n1039) );
  XOR2xp5r_ASAP7_6t_L U379 ( .A(n124), .B(n126), .Y(n64) );
  XOR2xp5r_ASAP7_6t_L U380 ( .A(n127), .B(n128), .Y(n63) );
  INVx1_ASAP7_6t_L U381 ( .A(n129), .Y(n127) );
  INVx1_ASAP7_6t_L U382 ( .A(n126), .Y(n125) );
  XOR2xp5r_ASAP7_6t_L U383 ( .A(n121), .B(n120), .Y(n126) );
  XOR2xp5r_ASAP7_6t_L U384 ( .A(n122), .B(n123), .Y(n120) );
  AO22x1_ASAP7_6t_L U385 ( .A1(n130), .A2(n131), .B1(n103), .B2(n104), .Y(n123) );
  XOR2xp5r_ASAP7_6t_L U386 ( .A(n131), .B(n130), .Y(n104) );
  XOR2xp5r_ASAP7_6t_L U387 ( .A(n132), .B(n133), .Y(n103) );
  XOR2xp5r_ASAP7_6t_L U388 ( .A(n134), .B(n135), .Y(n131) );
  XOR2xp5r_ASAP7_6t_L U389 ( .A(n136), .B(n137), .Y(n130) );
  OAI22xp5_ASAP7_6t_L U390 ( .A1(n138), .A2(n139), .B1(n140), .B2(n141), .Y(
        n122) );
  INVx1_ASAP7_6t_L U391 ( .A(n142), .Y(n138) );
  XOR2xp5r_ASAP7_6t_L U392 ( .A(n143), .B(n144), .Y(n121) );
  AOI22xp25_ASAP7_6t_L U393 ( .A1(n145), .A2(n146), .B1(n107), .B2(n106), .Y(
        n124) );
  XOR2xp5r_ASAP7_6t_L U394 ( .A(n140), .B(n141), .Y(n106) );
  XOR2xp5r_ASAP7_6t_L U395 ( .A(n142), .B(n139), .Y(n141) );
  AOI22xp25_ASAP7_6t_L U396 ( .A1(n147), .A2(n148), .B1(n149), .B2(n150), .Y(
        n139) );
  OAI22xp5_ASAP7_6t_L U397 ( .A1(n151), .A2(n152), .B1(n153), .B2(n154), .Y(
        n142) );
  AOI22xp25_ASAP7_6t_L U398 ( .A1(n155), .A2(n156), .B1(n157), .B2(n158), .Y(
        n140) );
  XOR2xp5r_ASAP7_6t_L U399 ( .A(n145), .B(n146), .Y(n107) );
  AO22x1_ASAP7_6t_L U400 ( .A1(n159), .A2(n160), .B1(n161), .B2(n162), .Y(n146) );
  AO22x1_ASAP7_6t_L U401 ( .A1(n163), .A2(n164), .B1(n165), .B2(n166), .Y(n145) );
  OAI22xp5_ASAP7_6t_L U402 ( .A1(n167), .A2(n168), .B1(n59), .B2(n60), .Y(
        n1040) );
  XOR2xp5r_ASAP7_6t_L U403 ( .A(n169), .B(n167), .Y(n60) );
  XOR2xp5r_ASAP7_6t_L U404 ( .A(n170), .B(n171), .Y(n59) );
  INVx1_ASAP7_6t_L U405 ( .A(n172), .Y(n170) );
  INVx1_ASAP7_6t_L U406 ( .A(n169), .Y(n168) );
  XOR2xp5r_ASAP7_6t_L U407 ( .A(n173), .B(n174), .Y(n169) );
  AOI22xp25_ASAP7_6t_L U408 ( .A1(n175), .A2(n176), .B1(n118), .B2(n119), .Y(
        n167) );
  XOR2xp5r_ASAP7_6t_L U409 ( .A(n177), .B(n178), .Y(n119) );
  XOR2xp5r_ASAP7_6t_L U410 ( .A(n175), .B(n176), .Y(n118) );
  AO22x1_ASAP7_6t_L U411 ( .A1(n179), .A2(n180), .B1(n129), .B2(n128), .Y(n176) );
  XOR2xp5r_ASAP7_6t_L U412 ( .A(n180), .B(n179), .Y(n128) );
  XOR2xp5r_ASAP7_6t_L U413 ( .A(n181), .B(n182), .Y(n129) );
  XOR2xp5r_ASAP7_6t_L U414 ( .A(n183), .B(n184), .Y(n180) );
  XOR2xp5r_ASAP7_6t_L U415 ( .A(n185), .B(n186), .Y(n179) );
  OAI22xp5_ASAP7_6t_L U416 ( .A1(n187), .A2(n188), .B1(n143), .B2(n144), .Y(
        n175) );
  XOR2xp5r_ASAP7_6t_L U417 ( .A(n189), .B(n188), .Y(n144) );
  INVx1_ASAP7_6t_L U418 ( .A(n187), .Y(n189) );
  AOI22xp25_ASAP7_6t_L U419 ( .A1(n190), .A2(n191), .B1(n132), .B2(n133), .Y(
        n143) );
  NOR2xp5_ASAP7_6t_L U420 ( .A(n90), .B(n41), .Y(n133) );
  XOR2xp5r_ASAP7_6t_L U421 ( .A(n190), .B(n191), .Y(n132) );
  XOR2xp5r_ASAP7_6t_L U422 ( .A(n192), .B(n193), .Y(n191) );
  XOR2xp5r_ASAP7_6t_L U423 ( .A(n194), .B(n195), .Y(n190) );
  AOI22xp25_ASAP7_6t_L U424 ( .A1(n196), .A2(n197), .B1(n136), .B2(n137), .Y(
        n188) );
  XOR2xp5r_ASAP7_6t_L U425 ( .A(n196), .B(n197), .Y(n137) );
  XOR2xp5r_ASAP7_6t_L U426 ( .A(n198), .B(n199), .Y(n136) );
  XOR2xp5r_ASAP7_6t_L U427 ( .A(n200), .B(n201), .Y(n197) );
  OAI22xp5_ASAP7_6t_L U428 ( .A1(n202), .A2(n203), .B1(n204), .B2(n205), .Y(
        n196) );
  AOI22xp25_ASAP7_6t_L U429 ( .A1(n206), .A2(n207), .B1(n134), .B2(n135), .Y(
        n187) );
  XOR2xp5r_ASAP7_6t_L U430 ( .A(n207), .B(n206), .Y(n135) );
  OAI22xp5_ASAP7_6t_L U431 ( .A1(n208), .A2(n209), .B1(n210), .B2(n211), .Y(
        n134) );
  OAI22xp5_ASAP7_6t_L U432 ( .A1(n212), .A2(n213), .B1(n214), .B2(n215), .Y(
        n207) );
  OAI22xp5_ASAP7_6t_L U433 ( .A1(n216), .A2(n217), .B1(n218), .B2(n219), .Y(
        n206) );
  INVx1_ASAP7_6t_L U434 ( .A(n220), .Y(n219) );
  OAI22xp5_ASAP7_6t_L U435 ( .A1(n221), .A2(n222), .B1(n58), .B2(n57), .Y(
        n1041) );
  INVx1_ASAP7_6t_L U436 ( .A(n223), .Y(n57) );
  XOR2xp5r_ASAP7_6t_L U437 ( .A(n224), .B(n225), .Y(n223) );
  XOR2xp5r_ASAP7_6t_L U438 ( .A(n226), .B(n221), .Y(n58) );
  INVx1_ASAP7_6t_L U439 ( .A(n226), .Y(n222) );
  XOR2xp5r_ASAP7_6t_L U440 ( .A(n227), .B(n228), .Y(n226) );
  OA22x1_ASAP7_6t_L U441 ( .A1(n229), .A2(n230), .B1(n174), .B2(n173), .Y(n221) );
  XOR2xp5r_ASAP7_6t_L U442 ( .A(n231), .B(n232), .Y(n173) );
  XOR2xp5r_ASAP7_6t_L U443 ( .A(n233), .B(n230), .Y(n174) );
  INVx1_ASAP7_6t_L U444 ( .A(n229), .Y(n233) );
  AOI22xp25_ASAP7_6t_L U445 ( .A1(n234), .A2(n235), .B1(n117), .B2(n116), .Y(
        n230) );
  XOR2xp5r_ASAP7_6t_L U446 ( .A(n234), .B(n235), .Y(n116) );
  XOR2xp5r_ASAP7_6t_L U447 ( .A(n236), .B(n237), .Y(n117) );
  XOR2xp5r_ASAP7_6t_L U448 ( .A(n238), .B(n239), .Y(n235) );
  XOR2xp5r_ASAP7_6t_L U449 ( .A(n240), .B(n241), .Y(n234) );
  AOI22xp25_ASAP7_6t_L U450 ( .A1(n242), .A2(n243), .B1(n178), .B2(n177), .Y(
        n229) );
  XOR2xp5r_ASAP7_6t_L U451 ( .A(n242), .B(n243), .Y(n177) );
  OAI22xp5_ASAP7_6t_L U452 ( .A1(n244), .A2(n245), .B1(n181), .B2(n182), .Y(
        n178) );
  NAND2xp5R_ASAP7_6t_L U453 ( .A(b[1]), .B(a[15]), .Y(n182) );
  XOR2xp5r_ASAP7_6t_L U454 ( .A(n246), .B(n245), .Y(n181) );
  XOR2xp5r_ASAP7_6t_L U455 ( .A(n247), .B(n248), .Y(n245) );
  INVx1_ASAP7_6t_L U456 ( .A(n246), .Y(n244) );
  XOR2xp5r_ASAP7_6t_L U457 ( .A(n249), .B(n250), .Y(n246) );
  AO22x1_ASAP7_6t_L U458 ( .A1(n251), .A2(n252), .B1(n185), .B2(n186), .Y(n243) );
  XOR2xp5r_ASAP7_6t_L U459 ( .A(n251), .B(n252), .Y(n186) );
  XOR2xp5r_ASAP7_6t_L U460 ( .A(n253), .B(n254), .Y(n185) );
  XOR2xp5r_ASAP7_6t_L U461 ( .A(n255), .B(n256), .Y(n252) );
  OAI22xp5_ASAP7_6t_L U462 ( .A1(n257), .A2(n258), .B1(n192), .B2(n193), .Y(
        n251) );
  NAND2xp5R_ASAP7_6t_L U463 ( .A(b[1]), .B(a[14]), .Y(n193) );
  INVx1_ASAP7_6t_L U464 ( .A(n259), .Y(n192) );
  XOR2xp5r_ASAP7_6t_L U465 ( .A(n257), .B(n258), .Y(n259) );
  NAND2xp5R_ASAP7_6t_L U466 ( .A(b[3]), .B(a[12]), .Y(n258) );
  NAND2xp5R_ASAP7_6t_L U467 ( .A(b[2]), .B(a[13]), .Y(n257) );
  AO22x1_ASAP7_6t_L U468 ( .A1(n260), .A2(n261), .B1(n183), .B2(n184), .Y(n242) );
  XOR2xp5r_ASAP7_6t_L U469 ( .A(n261), .B(n260), .Y(n184) );
  AO22x1_ASAP7_6t_L U470 ( .A1(n262), .A2(n263), .B1(n194), .B2(n195), .Y(n183) );
  AND2x2_ASAP7_6t_L U471 ( .A(b[4]), .B(a[11]), .Y(n195) );
  XOR2xp5r_ASAP7_6t_L U472 ( .A(n262), .B(n263), .Y(n194) );
  AND2x2_ASAP7_6t_L U473 ( .A(b[6]), .B(a[9]), .Y(n263) );
  NOR2xp5_ASAP7_6t_L U474 ( .A(n264), .B(n265), .Y(n262) );
  OAI22xp5_ASAP7_6t_L U475 ( .A1(n266), .A2(n267), .B1(n199), .B2(n198), .Y(
        n261) );
  NAND2xp5R_ASAP7_6t_L U476 ( .A(b[7]), .B(a[8]), .Y(n198) );
  XOR2xp5r_ASAP7_6t_L U477 ( .A(n267), .B(n268), .Y(n199) );
  XOR2xp5r_ASAP7_6t_L U478 ( .A(n269), .B(n270), .Y(n267) );
  NOR2xp5_ASAP7_6t_L U479 ( .A(n271), .B(n272), .Y(n269) );
  INVx1_ASAP7_6t_L U480 ( .A(n268), .Y(n266) );
  XOR2xp5r_ASAP7_6t_L U481 ( .A(n273), .B(n274), .Y(n268) );
  OAI22xp5_ASAP7_6t_L U482 ( .A1(n275), .A2(n276), .B1(n201), .B2(n200), .Y(
        n260) );
  XOR2xp5r_ASAP7_6t_L U483 ( .A(n275), .B(n277), .Y(n200) );
  XOR2xp5r_ASAP7_6t_L U484 ( .A(n278), .B(n279), .Y(n201) );
  INVx1_ASAP7_6t_L U485 ( .A(n277), .Y(n276) );
  NOR3x1f_ASAP7_6t_L U486 ( .A(n280), .B(n281), .C(n89), .Y(n277) );
  AOI22xp25_ASAP7_6t_L U487 ( .A1(n282), .A2(n283), .B1(n284), .B2(n285), .Y(
        n275) );
  OAI22xp5_ASAP7_6t_L U488 ( .A1(n286), .A2(n287), .B1(n55), .B2(n56), .Y(
        n1042) );
  XOR2xp5r_ASAP7_6t_L U489 ( .A(n288), .B(n286), .Y(n56) );
  INVx1_ASAP7_6t_L U490 ( .A(n287), .Y(n288) );
  XOR2xp5r_ASAP7_6t_L U491 ( .A(n289), .B(n290), .Y(n55) );
  INVx1_ASAP7_6t_L U492 ( .A(n291), .Y(n289) );
  XOR2xp5r_ASAP7_6t_L U493 ( .A(n292), .B(n293), .Y(n287) );
  AOI22xp25_ASAP7_6t_L U494 ( .A1(n294), .A2(n295), .B1(n228), .B2(n227), .Y(
        n286) );
  XOR2xp5r_ASAP7_6t_L U495 ( .A(n296), .B(n297), .Y(n227) );
  XOR2xp5r_ASAP7_6t_L U496 ( .A(n294), .B(n295), .Y(n228) );
  AO22x1_ASAP7_6t_L U497 ( .A1(n298), .A2(n299), .B1(n172), .B2(n171), .Y(n295) );
  XOR2xp5r_ASAP7_6t_L U498 ( .A(n298), .B(n299), .Y(n171) );
  XOR2xp5r_ASAP7_6t_L U499 ( .A(n300), .B(n301), .Y(n172) );
  XOR2xp5r_ASAP7_6t_L U500 ( .A(n302), .B(n303), .Y(n299) );
  XOR2xp5r_ASAP7_6t_L U501 ( .A(n304), .B(n305), .Y(n298) );
  OAI22xp5_ASAP7_6t_L U502 ( .A1(n306), .A2(n307), .B1(n308), .B2(n231), .Y(
        n294) );
  XOR2xp5r_ASAP7_6t_L U503 ( .A(n307), .B(n309), .Y(n231) );
  INVx1_ASAP7_6t_L U504 ( .A(n232), .Y(n308) );
  OAI22xp5_ASAP7_6t_L U505 ( .A1(n310), .A2(n311), .B1(n236), .B2(n237), .Y(
        n232) );
  NAND2xp5R_ASAP7_6t_L U506 ( .A(b[2]), .B(a[15]), .Y(n237) );
  XOR2xp5r_ASAP7_6t_L U507 ( .A(n312), .B(n311), .Y(n236) );
  INVx1_ASAP7_6t_L U508 ( .A(n310), .Y(n312) );
  XOR2xp5r_ASAP7_6t_L U509 ( .A(n313), .B(n314), .Y(n311) );
  XOR2xp5r_ASAP7_6t_L U510 ( .A(n315), .B(n316), .Y(n310) );
  AOI22xp25_ASAP7_6t_L U511 ( .A1(n317), .A2(n318), .B1(n240), .B2(n241), .Y(
        n307) );
  XOR2xp5r_ASAP7_6t_L U512 ( .A(n317), .B(n318), .Y(n241) );
  XOR2xp5r_ASAP7_6t_L U513 ( .A(n319), .B(n320), .Y(n240) );
  XOR2xp5r_ASAP7_6t_L U514 ( .A(n321), .B(n322), .Y(n318) );
  OAI22xp5_ASAP7_6t_L U515 ( .A1(n323), .A2(n324), .B1(n325), .B2(n248), .Y(
        n317) );
  NAND2xp5R_ASAP7_6t_L U516 ( .A(b[2]), .B(a[14]), .Y(n248) );
  INVx1_ASAP7_6t_L U517 ( .A(n247), .Y(n325) );
  XOR2xp5r_ASAP7_6t_L U518 ( .A(n324), .B(n323), .Y(n247) );
  NAND2xp5R_ASAP7_6t_L U519 ( .A(b[4]), .B(a[12]), .Y(n324) );
  NAND2xp5R_ASAP7_6t_L U520 ( .A(b[3]), .B(a[13]), .Y(n323) );
  INVx1_ASAP7_6t_L U521 ( .A(n309), .Y(n306) );
  OAI22xp5_ASAP7_6t_L U522 ( .A1(n326), .A2(n327), .B1(n238), .B2(n239), .Y(
        n309) );
  XOR2xp5r_ASAP7_6t_L U523 ( .A(n328), .B(n326), .Y(n239) );
  INVx1_ASAP7_6t_L U524 ( .A(n327), .Y(n328) );
  AOI22xp25_ASAP7_6t_L U525 ( .A1(n329), .A2(n330), .B1(n249), .B2(n250), .Y(
        n238) );
  AND2x2_ASAP7_6t_L U526 ( .A(b[5]), .B(a[11]), .Y(n250) );
  XOR2xp5r_ASAP7_6t_L U527 ( .A(n329), .B(n330), .Y(n249) );
  AND2x2_ASAP7_6t_L U528 ( .A(b[7]), .B(a[9]), .Y(n330) );
  NOR2xp5_ASAP7_6t_L U529 ( .A(n331), .B(n265), .Y(n329) );
  AOI22xp25_ASAP7_6t_L U530 ( .A1(n332), .A2(n333), .B1(n254), .B2(n253), .Y(
        n327) );
  XOR2xp5r_ASAP7_6t_L U531 ( .A(n332), .B(n333), .Y(n253) );
  XOR2xp5r_ASAP7_6t_L U532 ( .A(n334), .B(n335), .Y(n254) );
  NAND2xp5R_ASAP7_6t_L U533 ( .A(b[8]), .B(a[8]), .Y(n334) );
  XOR2xp5r_ASAP7_6t_L U534 ( .A(n336), .B(n337), .Y(n333) );
  XOR2xp5r_ASAP7_6t_L U535 ( .A(n338), .B(n339), .Y(n332) );
  AOI22xp25_ASAP7_6t_L U536 ( .A1(n340), .A2(n341), .B1(n255), .B2(n256), .Y(
        n326) );
  NOR3x1f_ASAP7_6t_L U537 ( .A(n270), .B(n271), .C(n272), .Y(n256) );
  NAND2xp5R_ASAP7_6t_L U538 ( .A(a[6]), .B(b[9]), .Y(n270) );
  XOR2xp5r_ASAP7_6t_L U539 ( .A(n341), .B(n340), .Y(n255) );
  AO22x1_ASAP7_6t_L U540 ( .A1(n342), .A2(n343), .B1(n273), .B2(n274), .Y(n341) );
  NOR2xp5_ASAP7_6t_L U541 ( .A(n344), .B(n281), .Y(n274) );
  XOR2xp5r_ASAP7_6t_L U542 ( .A(n343), .B(n342), .Y(n273) );
  NOR2xp5_ASAP7_6t_L U543 ( .A(n345), .B(n42), .Y(n343) );
  AND2x2_ASAP7_6t_L U544 ( .A(a[4]), .B(b[11]), .Y(n342) );
  OAI22xp5_ASAP7_6t_L U545 ( .A1(n346), .A2(n347), .B1(n348), .B2(n279), .Y(
        n340) );
  NAND2xp5R_ASAP7_6t_L U546 ( .A(a[2]), .B(b[13]), .Y(n279) );
  INVx1_ASAP7_6t_L U547 ( .A(n278), .Y(n348) );
  XOR2xp5r_ASAP7_6t_L U548 ( .A(n347), .B(n346), .Y(n278) );
  NAND2xp5R_ASAP7_6t_L U549 ( .A(a[0]), .B(b[15]), .Y(n347) );
  NAND2xp5R_ASAP7_6t_L U550 ( .A(a[1]), .B(b[14]), .Y(n346) );
  OAI22xp5_ASAP7_6t_L U551 ( .A1(n349), .A2(n350), .B1(n54), .B2(n53), .Y(
        n1043) );
  INVx1_ASAP7_6t_L U552 ( .A(n351), .Y(n53) );
  XOR2xp5r_ASAP7_6t_L U553 ( .A(n352), .B(n353), .Y(n351) );
  XOR2xp5r_ASAP7_6t_L U554 ( .A(n354), .B(n349), .Y(n54) );
  INVx1_ASAP7_6t_L U555 ( .A(n354), .Y(n350) );
  XOR2xp5r_ASAP7_6t_L U556 ( .A(n355), .B(n356), .Y(n354) );
  OA22x1_ASAP7_6t_L U557 ( .A1(n357), .A2(n358), .B1(n359), .B2(n292), .Y(n349) );
  XOR2xp5r_ASAP7_6t_L U558 ( .A(n360), .B(n361), .Y(n292) );
  INVx1_ASAP7_6t_L U559 ( .A(n293), .Y(n359) );
  XOR2xp5r_ASAP7_6t_L U560 ( .A(n357), .B(n358), .Y(n293) );
  AOI22xp25_ASAP7_6t_L U561 ( .A1(n362), .A2(n363), .B1(n224), .B2(n225), .Y(
        n358) );
  XOR2xp5r_ASAP7_6t_L U562 ( .A(n362), .B(n363), .Y(n225) );
  XOR2xp5r_ASAP7_6t_L U563 ( .A(n364), .B(n365), .Y(n224) );
  XOR2xp5r_ASAP7_6t_L U564 ( .A(n366), .B(n367), .Y(n363) );
  XOR2xp5r_ASAP7_6t_L U565 ( .A(n368), .B(n369), .Y(n362) );
  AOI22xp25_ASAP7_6t_L U566 ( .A1(n370), .A2(n371), .B1(n297), .B2(n296), .Y(
        n357) );
  XOR2xp5r_ASAP7_6t_L U567 ( .A(n371), .B(n370), .Y(n296) );
  OAI22xp5_ASAP7_6t_L U568 ( .A1(n372), .A2(n373), .B1(n300), .B2(n301), .Y(
        n297) );
  NAND2xp5R_ASAP7_6t_L U569 ( .A(b[3]), .B(a[15]), .Y(n301) );
  XOR2xp5r_ASAP7_6t_L U570 ( .A(n374), .B(n373), .Y(n300) );
  XOR2xp5r_ASAP7_6t_L U571 ( .A(n375), .B(n376), .Y(n373) );
  INVx1_ASAP7_6t_L U572 ( .A(n374), .Y(n372) );
  XOR2xp5r_ASAP7_6t_L U573 ( .A(n377), .B(n378), .Y(n374) );
  AO22x1_ASAP7_6t_L U574 ( .A1(n379), .A2(n380), .B1(n304), .B2(n305), .Y(n371) );
  XOR2xp5r_ASAP7_6t_L U575 ( .A(n379), .B(n380), .Y(n305) );
  XOR2xp5r_ASAP7_6t_L U576 ( .A(n381), .B(n382), .Y(n304) );
  XOR2xp5r_ASAP7_6t_L U577 ( .A(n383), .B(n384), .Y(n380) );
  OAI22xp5_ASAP7_6t_L U578 ( .A1(n385), .A2(n386), .B1(n387), .B2(n314), .Y(
        n379) );
  NAND2xp5R_ASAP7_6t_L U579 ( .A(b[3]), .B(a[14]), .Y(n314) );
  INVx1_ASAP7_6t_L U580 ( .A(n313), .Y(n387) );
  XOR2xp5r_ASAP7_6t_L U581 ( .A(n385), .B(n386), .Y(n313) );
  NAND2xp5R_ASAP7_6t_L U582 ( .A(b[5]), .B(a[12]), .Y(n386) );
  NAND2xp5R_ASAP7_6t_L U583 ( .A(b[4]), .B(a[13]), .Y(n385) );
  OAI22xp5_ASAP7_6t_L U584 ( .A1(n388), .A2(n389), .B1(n302), .B2(n303), .Y(
        n370) );
  INVx1_ASAP7_6t_L U585 ( .A(n390), .Y(n303) );
  XOR2xp5r_ASAP7_6t_L U586 ( .A(n389), .B(n388), .Y(n390) );
  OA22x1_ASAP7_6t_L U587 ( .A1(n391), .A2(n392), .B1(n393), .B2(n316), .Y(n302) );
  NAND2xp5R_ASAP7_6t_L U588 ( .A(b[6]), .B(a[11]), .Y(n316) );
  INVx1_ASAP7_6t_L U589 ( .A(n315), .Y(n393) );
  XOR2xp5r_ASAP7_6t_L U590 ( .A(n391), .B(n392), .Y(n315) );
  NAND2xp5R_ASAP7_6t_L U591 ( .A(b[8]), .B(a[9]), .Y(n392) );
  NAND2xp5R_ASAP7_6t_L U592 ( .A(b[7]), .B(a[10]), .Y(n391) );
  AOI22xp25_ASAP7_6t_L U593 ( .A1(n394), .A2(n395), .B1(n319), .B2(n320), .Y(
        n389) );
  AND2x2_ASAP7_6t_L U594 ( .A(a[8]), .B(b[9]), .Y(n320) );
  XOR2xp5r_ASAP7_6t_L U595 ( .A(n395), .B(n394), .Y(n319) );
  XOR2xp5r_ASAP7_6t_L U596 ( .A(n396), .B(n397), .Y(n395) );
  XOR2xp5r_ASAP7_6t_L U597 ( .A(n398), .B(n399), .Y(n394) );
  AOI22xp25_ASAP7_6t_L U598 ( .A1(n400), .A2(n401), .B1(n321), .B2(n322), .Y(
        n388) );
  NOR3x1f_ASAP7_6t_L U599 ( .A(n335), .B(n271), .C(n402), .Y(n322) );
  NAND2xp5R_ASAP7_6t_L U600 ( .A(a[7]), .B(b[9]), .Y(n335) );
  XOR2xp5r_ASAP7_6t_L U601 ( .A(n401), .B(n400), .Y(n321) );
  OAI22xp5_ASAP7_6t_L U602 ( .A1(n403), .A2(n404), .B1(n336), .B2(n337), .Y(
        n401) );
  NAND2xp5R_ASAP7_6t_L U603 ( .A(a[6]), .B(b[10]), .Y(n337) );
  INVx1_ASAP7_6t_L U604 ( .A(n405), .Y(n336) );
  XOR2xp5r_ASAP7_6t_L U605 ( .A(n403), .B(n404), .Y(n405) );
  NAND2xp5R_ASAP7_6t_L U606 ( .A(a[4]), .B(b[12]), .Y(n404) );
  NAND2xp5R_ASAP7_6t_L U607 ( .A(a[5]), .B(b[11]), .Y(n403) );
  OAI22xp5_ASAP7_6t_L U608 ( .A1(n406), .A2(n407), .B1(n338), .B2(n339), .Y(
        n400) );
  NAND2xp5R_ASAP7_6t_L U609 ( .A(a[3]), .B(b[13]), .Y(n339) );
  XOR2xp5r_ASAP7_6t_L U610 ( .A(n408), .B(n407), .Y(n338) );
  NAND2xp5R_ASAP7_6t_L U611 ( .A(a[1]), .B(b[15]), .Y(n407) );
  INVx1_ASAP7_6t_L U612 ( .A(n408), .Y(n406) );
  NOR2xp5_ASAP7_6t_L U613 ( .A(n95), .B(n409), .Y(n408) );
  OAI22xp5_ASAP7_6t_L U614 ( .A1(n410), .A2(n411), .B1(n51), .B2(n52), .Y(
        n1044) );
  XOR2xp5r_ASAP7_6t_L U615 ( .A(n412), .B(n410), .Y(n52) );
  XOR2xp5r_ASAP7_6t_L U616 ( .A(n413), .B(n414), .Y(n51) );
  INVx1_ASAP7_6t_L U617 ( .A(n412), .Y(n411) );
  XOR2xp5r_ASAP7_6t_L U618 ( .A(n415), .B(n416), .Y(n412) );
  AOI22xp25_ASAP7_6t_L U619 ( .A1(n417), .A2(n418), .B1(n355), .B2(n356), .Y(
        n410) );
  XOR2xp5r_ASAP7_6t_L U620 ( .A(n419), .B(n420), .Y(n356) );
  XOR2xp5r_ASAP7_6t_L U621 ( .A(n418), .B(n417), .Y(n355) );
  AO22x1_ASAP7_6t_L U622 ( .A1(n421), .A2(n422), .B1(n291), .B2(n290), .Y(n418) );
  XOR2xp5r_ASAP7_6t_L U623 ( .A(n421), .B(n422), .Y(n290) );
  XOR2xp5r_ASAP7_6t_L U624 ( .A(n423), .B(n424), .Y(n291) );
  XOR2xp5r_ASAP7_6t_L U625 ( .A(n425), .B(n426), .Y(n422) );
  XOR2xp5r_ASAP7_6t_L U626 ( .A(n427), .B(n428), .Y(n421) );
  OAI22xp5_ASAP7_6t_L U627 ( .A1(n429), .A2(n430), .B1(n361), .B2(n431), .Y(
        n417) );
  INVx1_ASAP7_6t_L U628 ( .A(n360), .Y(n431) );
  XOR2xp5r_ASAP7_6t_L U629 ( .A(n430), .B(n429), .Y(n360) );
  OA22x1_ASAP7_6t_L U630 ( .A1(n432), .A2(n433), .B1(n364), .B2(n365), .Y(n361) );
  NAND2xp5R_ASAP7_6t_L U631 ( .A(b[4]), .B(a[15]), .Y(n365) );
  XOR2xp5r_ASAP7_6t_L U632 ( .A(n434), .B(n432), .Y(n364) );
  INVx1_ASAP7_6t_L U633 ( .A(n434), .Y(n433) );
  XOR2xp5r_ASAP7_6t_L U634 ( .A(n435), .B(n436), .Y(n434) );
  XOR2xp5r_ASAP7_6t_L U635 ( .A(n437), .B(n438), .Y(n432) );
  AOI22xp25_ASAP7_6t_L U636 ( .A1(n439), .A2(n440), .B1(n368), .B2(n369), .Y(
        n430) );
  XOR2xp5r_ASAP7_6t_L U637 ( .A(n439), .B(n440), .Y(n369) );
  XOR2xp5r_ASAP7_6t_L U638 ( .A(n441), .B(n442), .Y(n368) );
  XOR2xp5r_ASAP7_6t_L U639 ( .A(n443), .B(n444), .Y(n440) );
  OAI22xp5_ASAP7_6t_L U640 ( .A1(n445), .A2(n446), .B1(n447), .B2(n376), .Y(
        n439) );
  NAND2xp5R_ASAP7_6t_L U641 ( .A(b[4]), .B(a[14]), .Y(n376) );
  INVx1_ASAP7_6t_L U642 ( .A(n375), .Y(n447) );
  XOR2xp5r_ASAP7_6t_L U643 ( .A(n445), .B(n446), .Y(n375) );
  NAND2xp5R_ASAP7_6t_L U644 ( .A(b[6]), .B(a[12]), .Y(n446) );
  NAND2xp5R_ASAP7_6t_L U645 ( .A(b[5]), .B(a[13]), .Y(n445) );
  AOI22xp25_ASAP7_6t_L U646 ( .A1(n448), .A2(n449), .B1(n366), .B2(n367), .Y(
        n429) );
  XOR2xp5r_ASAP7_6t_L U647 ( .A(n449), .B(n448), .Y(n367) );
  OAI22xp5_ASAP7_6t_L U648 ( .A1(n450), .A2(n451), .B1(n377), .B2(n378), .Y(
        n366) );
  NAND2xp5R_ASAP7_6t_L U649 ( .A(b[7]), .B(a[11]), .Y(n378) );
  INVx1_ASAP7_6t_L U650 ( .A(n452), .Y(n377) );
  XOR2xp5r_ASAP7_6t_L U651 ( .A(n451), .B(n450), .Y(n452) );
  NAND2xp5R_ASAP7_6t_L U652 ( .A(b[9]), .B(a[9]), .Y(n451) );
  NAND2xp5R_ASAP7_6t_L U653 ( .A(b[8]), .B(a[10]), .Y(n450) );
  OAI22xp5_ASAP7_6t_L U654 ( .A1(n453), .A2(n454), .B1(n381), .B2(n382), .Y(
        n449) );
  NAND2xp5R_ASAP7_6t_L U655 ( .A(a[8]), .B(b[10]), .Y(n382) );
  XOR2xp5r_ASAP7_6t_L U656 ( .A(n455), .B(n454), .Y(n381) );
  INVx1_ASAP7_6t_L U657 ( .A(n453), .Y(n455) );
  NAND2xp5R_ASAP7_6t_L U658 ( .A(a[6]), .B(b[12]), .Y(n454) );
  NAND2xp5R_ASAP7_6t_L U659 ( .A(a[7]), .B(b[11]), .Y(n453) );
  AO22x1_ASAP7_6t_L U660 ( .A1(n456), .A2(n457), .B1(n384), .B2(n383), .Y(n448) );
  XOR2xp5r_ASAP7_6t_L U661 ( .A(n457), .B(n456), .Y(n383) );
  XOR2xp5r_ASAP7_6t_L U662 ( .A(n458), .B(n459), .Y(n384) );
  OAI22xp5_ASAP7_6t_L U663 ( .A1(n460), .A2(n461), .B1(n396), .B2(n397), .Y(
        n457) );
  NAND2xp5R_ASAP7_6t_L U664 ( .A(a[7]), .B(b[10]), .Y(n397) );
  XOR2xp5r_ASAP7_6t_L U665 ( .A(n462), .B(n461), .Y(n396) );
  INVx1_ASAP7_6t_L U666 ( .A(n460), .Y(n462) );
  NAND2xp5R_ASAP7_6t_L U667 ( .A(a[5]), .B(b[12]), .Y(n461) );
  NAND2xp5R_ASAP7_6t_L U668 ( .A(a[6]), .B(b[11]), .Y(n460) );
  OAI22xp5_ASAP7_6t_L U669 ( .A1(n463), .A2(n464), .B1(n398), .B2(n399), .Y(
        n456) );
  NAND2xp5R_ASAP7_6t_L U670 ( .A(a[4]), .B(b[13]), .Y(n399) );
  XOR2xp5r_ASAP7_6t_L U671 ( .A(n465), .B(n464), .Y(n398) );
  INVx1_ASAP7_6t_L U672 ( .A(n463), .Y(n465) );
  NAND2xp5R_ASAP7_6t_L U673 ( .A(a[2]), .B(b[15]), .Y(n464) );
  NAND2xp5R_ASAP7_6t_L U674 ( .A(a[3]), .B(b[14]), .Y(n463) );
  OAI22xp5_ASAP7_6t_L U675 ( .A1(n466), .A2(n467), .B1(n50), .B2(n49), .Y(
        n1045) );
  INVx1_ASAP7_6t_L U676 ( .A(n468), .Y(n49) );
  XOR2xp5r_ASAP7_6t_L U677 ( .A(n469), .B(n470), .Y(n468) );
  XOR2xp5r_ASAP7_6t_L U678 ( .A(n471), .B(n466), .Y(n50) );
  INVx1_ASAP7_6t_L U679 ( .A(n471), .Y(n467) );
  XOR2xp5r_ASAP7_6t_L U680 ( .A(n472), .B(n473), .Y(n471) );
  AOI22xp25_ASAP7_6t_L U681 ( .A1(n474), .A2(n475), .B1(n416), .B2(n415), .Y(
        n466) );
  XOR2xp5r_ASAP7_6t_L U682 ( .A(n476), .B(n477), .Y(n415) );
  XOR2xp5r_ASAP7_6t_L U683 ( .A(n475), .B(n474), .Y(n416) );
  AO22x1_ASAP7_6t_L U684 ( .A1(n478), .A2(n479), .B1(n352), .B2(n353), .Y(n475) );
  XOR2xp5r_ASAP7_6t_L U685 ( .A(n478), .B(n479), .Y(n353) );
  XOR2xp5r_ASAP7_6t_L U686 ( .A(n480), .B(n481), .Y(n352) );
  XOR2xp5r_ASAP7_6t_L U687 ( .A(n482), .B(n483), .Y(n479) );
  XOR2xp5r_ASAP7_6t_L U688 ( .A(n484), .B(n485), .Y(n478) );
  OAI22xp5_ASAP7_6t_L U689 ( .A1(n486), .A2(n487), .B1(n419), .B2(n420), .Y(
        n474) );
  XOR2xp5r_ASAP7_6t_L U690 ( .A(n488), .B(n486), .Y(n420) );
  INVx1_ASAP7_6t_L U691 ( .A(n487), .Y(n488) );
  AOI22xp25_ASAP7_6t_L U692 ( .A1(n489), .A2(n490), .B1(n424), .B2(n423), .Y(
        n419) );
  NOR2xp5_ASAP7_6t_L U693 ( .A(n264), .B(n41), .Y(n423) );
  XOR2xp5r_ASAP7_6t_L U694 ( .A(n490), .B(n489), .Y(n424) );
  NOR2xp5_ASAP7_6t_L U695 ( .A(n331), .B(n491), .Y(n490) );
  XOR2xp5r_ASAP7_6t_L U696 ( .A(n492), .B(n493), .Y(n489) );
  AOI22xp25_ASAP7_6t_L U697 ( .A1(n494), .A2(n495), .B1(n427), .B2(n428), .Y(
        n487) );
  XOR2xp5r_ASAP7_6t_L U698 ( .A(n494), .B(n495), .Y(n428) );
  XOR2xp5r_ASAP7_6t_L U699 ( .A(n496), .B(n497), .Y(n427) );
  XOR2xp5r_ASAP7_6t_L U700 ( .A(n498), .B(n499), .Y(n495) );
  OAI22xp5_ASAP7_6t_L U701 ( .A1(n500), .A2(n501), .B1(n435), .B2(n436), .Y(
        n494) );
  NAND2xp5R_ASAP7_6t_L U702 ( .A(b[5]), .B(a[14]), .Y(n436) );
  XOR2xp5r_ASAP7_6t_L U703 ( .A(n502), .B(n501), .Y(n435) );
  INVx1_ASAP7_6t_L U704 ( .A(n500), .Y(n502) );
  NAND2xp5R_ASAP7_6t_L U705 ( .A(b[7]), .B(a[12]), .Y(n501) );
  NAND2xp5R_ASAP7_6t_L U706 ( .A(b[6]), .B(a[13]), .Y(n500) );
  AOI22xp25_ASAP7_6t_L U707 ( .A1(n503), .A2(n504), .B1(n425), .B2(n426), .Y(
        n486) );
  XOR2xp5r_ASAP7_6t_L U708 ( .A(n504), .B(n503), .Y(n426) );
  OAI22xp5_ASAP7_6t_L U709 ( .A1(n505), .A2(n506), .B1(n507), .B2(n438), .Y(
        n425) );
  NAND2xp5R_ASAP7_6t_L U710 ( .A(b[8]), .B(a[11]), .Y(n438) );
  INVx1_ASAP7_6t_L U711 ( .A(n437), .Y(n507) );
  XOR2xp5r_ASAP7_6t_L U712 ( .A(n505), .B(n506), .Y(n437) );
  NAND2xp5R_ASAP7_6t_L U713 ( .A(a[9]), .B(b[10]), .Y(n506) );
  NAND2xp5R_ASAP7_6t_L U714 ( .A(b[9]), .B(a[10]), .Y(n505) );
  OAI22xp5_ASAP7_6t_L U715 ( .A1(n508), .A2(n509), .B1(n441), .B2(n442), .Y(
        n504) );
  NAND2xp5R_ASAP7_6t_L U716 ( .A(a[8]), .B(b[11]), .Y(n442) );
  XOR2xp5r_ASAP7_6t_L U717 ( .A(n510), .B(n508), .Y(n441) );
  INVx1_ASAP7_6t_L U718 ( .A(n509), .Y(n510) );
  NAND2xp5R_ASAP7_6t_L U719 ( .A(a[6]), .B(b[13]), .Y(n509) );
  NAND2xp5R_ASAP7_6t_L U720 ( .A(a[7]), .B(b[12]), .Y(n508) );
  OAI22xp5_ASAP7_6t_L U721 ( .A1(n511), .A2(n512), .B1(n443), .B2(n444), .Y(
        n503) );
  NAND2xp5R_ASAP7_6t_L U722 ( .A(a[5]), .B(b[14]), .Y(n444) );
  XOR2xp5r_ASAP7_6t_L U723 ( .A(n513), .B(n512), .Y(n443) );
  INVx1_ASAP7_6t_L U724 ( .A(n511), .Y(n513) );
  NAND2xp5R_ASAP7_6t_L U725 ( .A(a[4]), .B(b[15]), .Y(n512) );
  AOI22xp25_ASAP7_6t_L U726 ( .A1(n514), .A2(n515), .B1(n458), .B2(n459), .Y(
        n511) );
  NOR2xp5_ASAP7_6t_L U727 ( .A(n344), .B(n516), .Y(n459) );
  XOR2xp5r_ASAP7_6t_L U728 ( .A(n515), .B(n514), .Y(n458) );
  NOR2xp5_ASAP7_6t_L U729 ( .A(n345), .B(n96), .Y(n515) );
  NOR2xp5_ASAP7_6t_L U730 ( .A(n89), .B(n409), .Y(n514) );
  OAI22xp5_ASAP7_6t_L U731 ( .A1(n517), .A2(n518), .B1(n47), .B2(n48), .Y(
        n1046) );
  XOR2xp5r_ASAP7_6t_L U732 ( .A(n519), .B(n517), .Y(n48) );
  XOR2xp5r_ASAP7_6t_L U733 ( .A(n520), .B(n521), .Y(n47) );
  INVx1_ASAP7_6t_L U734 ( .A(n522), .Y(n520) );
  INVx1_ASAP7_6t_L U735 ( .A(n519), .Y(n518) );
  XOR2xp5r_ASAP7_6t_L U736 ( .A(n523), .B(n524), .Y(n519) );
  AOI22xp25_ASAP7_6t_L U737 ( .A1(n525), .A2(n526), .B1(n472), .B2(n473), .Y(
        n517) );
  XOR2xp5r_ASAP7_6t_L U738 ( .A(n527), .B(n528), .Y(n473) );
  XOR2xp5r_ASAP7_6t_L U739 ( .A(n526), .B(n525), .Y(n472) );
  AO22x1_ASAP7_6t_L U740 ( .A1(n529), .A2(n530), .B1(n531), .B2(n414), .Y(n526) );
  XOR2xp5r_ASAP7_6t_L U741 ( .A(n530), .B(n529), .Y(n414) );
  INVx1_ASAP7_6t_L U742 ( .A(n413), .Y(n531) );
  XOR2xp5r_ASAP7_6t_L U743 ( .A(n532), .B(n533), .Y(n413) );
  XOR2xp5r_ASAP7_6t_L U744 ( .A(n534), .B(n535), .Y(n530) );
  XOR2xp5r_ASAP7_6t_L U745 ( .A(n536), .B(n537), .Y(n529) );
  OAI22xp5_ASAP7_6t_L U746 ( .A1(n538), .A2(n539), .B1(n476), .B2(n477), .Y(
        n525) );
  XOR2xp5r_ASAP7_6t_L U747 ( .A(n540), .B(n538), .Y(n477) );
  INVx1_ASAP7_6t_L U748 ( .A(n539), .Y(n540) );
  OA22x1_ASAP7_6t_L U749 ( .A1(n541), .A2(n542), .B1(n480), .B2(n481), .Y(n476) );
  NAND2xp5R_ASAP7_6t_L U750 ( .A(b[6]), .B(a[15]), .Y(n481) );
  XOR2xp5r_ASAP7_6t_L U751 ( .A(n543), .B(n542), .Y(n480) );
  INVx1_ASAP7_6t_L U752 ( .A(n541), .Y(n543) );
  NAND2xp5R_ASAP7_6t_L U753 ( .A(b[8]), .B(a[13]), .Y(n542) );
  NAND2xp5R_ASAP7_6t_L U754 ( .A(b[7]), .B(a[14]), .Y(n541) );
  AOI22xp25_ASAP7_6t_L U755 ( .A1(n544), .A2(n545), .B1(n484), .B2(n485), .Y(
        n539) );
  AND2x2_ASAP7_6t_L U756 ( .A(b[9]), .B(a[12]), .Y(n485) );
  XOR2xp5r_ASAP7_6t_L U757 ( .A(n544), .B(n545), .Y(n484) );
  XOR2xp5r_ASAP7_6t_L U758 ( .A(n546), .B(n547), .Y(n545) );
  XOR2xp5r_ASAP7_6t_L U759 ( .A(n548), .B(n549), .Y(n544) );
  AOI22xp25_ASAP7_6t_L U760 ( .A1(n550), .A2(n551), .B1(n483), .B2(n482), .Y(
        n538) );
  XOR2xp5r_ASAP7_6t_L U761 ( .A(n551), .B(n550), .Y(n482) );
  OAI22xp5_ASAP7_6t_L U762 ( .A1(n552), .A2(n553), .B1(n492), .B2(n493), .Y(
        n483) );
  NAND2xp5R_ASAP7_6t_L U763 ( .A(b[7]), .B(a[13]), .Y(n493) );
  INVx1_ASAP7_6t_L U764 ( .A(n554), .Y(n492) );
  XOR2xp5r_ASAP7_6t_L U765 ( .A(n553), .B(n552), .Y(n554) );
  NAND2xp5R_ASAP7_6t_L U766 ( .A(b[9]), .B(a[11]), .Y(n553) );
  NAND2xp5R_ASAP7_6t_L U767 ( .A(b[8]), .B(a[12]), .Y(n552) );
  OAI22xp5_ASAP7_6t_L U768 ( .A1(n555), .A2(n556), .B1(n496), .B2(n497), .Y(
        n551) );
  NAND2xp5R_ASAP7_6t_L U769 ( .A(b[10]), .B(a[10]), .Y(n497) );
  XOR2xp5r_ASAP7_6t_L U770 ( .A(n557), .B(n556), .Y(n496) );
  INVx1_ASAP7_6t_L U771 ( .A(n555), .Y(n557) );
  NAND2xp5R_ASAP7_6t_L U772 ( .A(a[8]), .B(b[12]), .Y(n556) );
  NAND2xp5R_ASAP7_6t_L U773 ( .A(a[9]), .B(b[11]), .Y(n555) );
  OAI22xp5_ASAP7_6t_L U774 ( .A1(n558), .A2(n559), .B1(n498), .B2(n499), .Y(
        n550) );
  NAND2xp5R_ASAP7_6t_L U775 ( .A(a[7]), .B(b[13]), .Y(n499) );
  INVx1_ASAP7_6t_L U776 ( .A(n560), .Y(n498) );
  XOR2xp5r_ASAP7_6t_L U777 ( .A(n558), .B(n559), .Y(n560) );
  NAND2xp5R_ASAP7_6t_L U778 ( .A(a[5]), .B(b[15]), .Y(n559) );
  NAND2xp5R_ASAP7_6t_L U779 ( .A(a[6]), .B(b[14]), .Y(n558) );
  OAI22xp5_ASAP7_6t_L U780 ( .A1(n561), .A2(n562), .B1(n45), .B2(n46), .Y(
        n1047) );
  XOR2xp5r_ASAP7_6t_L U781 ( .A(n563), .B(n561), .Y(n46) );
  XOR2xp5r_ASAP7_6t_L U782 ( .A(n564), .B(n565), .Y(n45) );
  INVx1_ASAP7_6t_L U783 ( .A(n563), .Y(n562) );
  XOR2xp5r_ASAP7_6t_L U784 ( .A(n566), .B(n567), .Y(n563) );
  AOI22xp25_ASAP7_6t_L U785 ( .A1(n568), .A2(n569), .B1(n523), .B2(n524), .Y(
        n561) );
  XOR2xp5r_ASAP7_6t_L U786 ( .A(n570), .B(n571), .Y(n524) );
  XOR2xp5r_ASAP7_6t_L U787 ( .A(n569), .B(n568), .Y(n523) );
  AO22x1_ASAP7_6t_L U788 ( .A1(n572), .A2(n573), .B1(n469), .B2(n470), .Y(n569) );
  XOR2xp5r_ASAP7_6t_L U789 ( .A(n572), .B(n573), .Y(n470) );
  XOR2xp5r_ASAP7_6t_L U790 ( .A(n574), .B(n575), .Y(n469) );
  XOR2xp5r_ASAP7_6t_L U791 ( .A(n576), .B(n577), .Y(n573) );
  XOR2xp5r_ASAP7_6t_L U792 ( .A(n578), .B(n579), .Y(n572) );
  AO22x1_ASAP7_6t_L U793 ( .A1(n580), .A2(n581), .B1(n527), .B2(n528), .Y(n568) );
  XOR2xp5r_ASAP7_6t_L U794 ( .A(n581), .B(n580), .Y(n528) );
  OAI22xp5_ASAP7_6t_L U795 ( .A1(n582), .A2(n583), .B1(n584), .B2(n533), .Y(
        n527) );
  NAND2xp5R_ASAP7_6t_L U796 ( .A(b[7]), .B(a[15]), .Y(n533) );
  INVx1_ASAP7_6t_L U797 ( .A(n532), .Y(n584) );
  XOR2xp5r_ASAP7_6t_L U798 ( .A(n583), .B(n582), .Y(n532) );
  NAND2xp5R_ASAP7_6t_L U799 ( .A(b[9]), .B(a[13]), .Y(n583) );
  NAND2xp5R_ASAP7_6t_L U800 ( .A(b[8]), .B(a[14]), .Y(n582) );
  OAI22xp5_ASAP7_6t_L U801 ( .A1(n585), .A2(n586), .B1(n534), .B2(n535), .Y(
        n581) );
  NAND2xp5R_ASAP7_6t_L U802 ( .A(b[10]), .B(a[12]), .Y(n535) );
  XOR2xp5r_ASAP7_6t_L U803 ( .A(n587), .B(n586), .Y(n534) );
  INVx1_ASAP7_6t_L U804 ( .A(n585), .Y(n587) );
  NAND2xp5R_ASAP7_6t_L U805 ( .A(a[10]), .B(b[12]), .Y(n586) );
  NAND2xp5R_ASAP7_6t_L U806 ( .A(a[11]), .B(b[11]), .Y(n585) );
  AO22x1_ASAP7_6t_L U807 ( .A1(n588), .A2(n589), .B1(n537), .B2(n536), .Y(n580) );
  XOR2xp5r_ASAP7_6t_L U808 ( .A(n589), .B(n588), .Y(n536) );
  XOR2xp5r_ASAP7_6t_L U809 ( .A(n590), .B(n591), .Y(n537) );
  OAI22xp5_ASAP7_6t_L U810 ( .A1(n592), .A2(n593), .B1(n546), .B2(n547), .Y(
        n589) );
  NAND2xp5R_ASAP7_6t_L U811 ( .A(b[10]), .B(a[11]), .Y(n547) );
  INVx1_ASAP7_6t_L U812 ( .A(n594), .Y(n546) );
  XOR2xp5r_ASAP7_6t_L U813 ( .A(n592), .B(n593), .Y(n594) );
  NAND2xp5R_ASAP7_6t_L U814 ( .A(a[9]), .B(b[12]), .Y(n593) );
  NAND2xp5R_ASAP7_6t_L U815 ( .A(a[10]), .B(b[11]), .Y(n592) );
  OAI22xp5_ASAP7_6t_L U816 ( .A1(n595), .A2(n596), .B1(n548), .B2(n549), .Y(
        n588) );
  NAND2xp5R_ASAP7_6t_L U817 ( .A(a[8]), .B(b[13]), .Y(n549) );
  XOR2xp5r_ASAP7_6t_L U818 ( .A(n597), .B(n595), .Y(n548) );
  INVx1_ASAP7_6t_L U819 ( .A(n596), .Y(n597) );
  NAND2xp5R_ASAP7_6t_L U820 ( .A(a[6]), .B(b[15]), .Y(n596) );
  NAND2xp5R_ASAP7_6t_L U821 ( .A(a[7]), .B(b[14]), .Y(n595) );
  OAI22xp5_ASAP7_6t_L U822 ( .A1(n598), .A2(n599), .B1(n43), .B2(n44), .Y(
        n1048) );
  XOR2xp5r_ASAP7_6t_L U823 ( .A(n600), .B(n598), .Y(n44) );
  XOR2xp5r_ASAP7_6t_L U824 ( .A(n601), .B(n602), .Y(n43) );
  INVx1_ASAP7_6t_L U825 ( .A(n600), .Y(n599) );
  XOR2xp5r_ASAP7_6t_L U826 ( .A(n603), .B(n604), .Y(n600) );
  AOI22xp25_ASAP7_6t_L U827 ( .A1(n605), .A2(n606), .B1(n566), .B2(n567), .Y(
        n598) );
  XOR2xp5r_ASAP7_6t_L U828 ( .A(n606), .B(n605), .Y(n567) );
  XOR2xp5r_ASAP7_6t_L U829 ( .A(n607), .B(n608), .Y(n566) );
  AO22x1_ASAP7_6t_L U830 ( .A1(n609), .A2(n610), .B1(n522), .B2(n521), .Y(n606) );
  AND2x2_ASAP7_6t_L U831 ( .A(b[9]), .B(a[15]), .Y(n521) );
  XOR2xp5r_ASAP7_6t_L U832 ( .A(n609), .B(n610), .Y(n522) );
  XOR2xp5r_ASAP7_6t_L U833 ( .A(n611), .B(n612), .Y(n610) );
  XOR2xp5r_ASAP7_6t_L U834 ( .A(n613), .B(n614), .Y(n609) );
  OAI22xp5_ASAP7_6t_L U835 ( .A1(n615), .A2(n616), .B1(n570), .B2(n571), .Y(
        n605) );
  XOR2xp5r_ASAP7_6t_L U836 ( .A(n616), .B(n617), .Y(n571) );
  OA22x1_ASAP7_6t_L U837 ( .A1(n618), .A2(n619), .B1(n574), .B2(n575), .Y(n570) );
  NAND2xp5R_ASAP7_6t_L U838 ( .A(b[8]), .B(a[15]), .Y(n575) );
  XOR2xp5r_ASAP7_6t_L U839 ( .A(n620), .B(n619), .Y(n574) );
  INVx1_ASAP7_6t_L U840 ( .A(n618), .Y(n620) );
  NAND2xp5R_ASAP7_6t_L U841 ( .A(b[10]), .B(a[13]), .Y(n619) );
  NAND2xp5R_ASAP7_6t_L U842 ( .A(b[9]), .B(a[14]), .Y(n618) );
  AOI22xp25_ASAP7_6t_L U843 ( .A1(n621), .A2(n622), .B1(n578), .B2(n579), .Y(
        n616) );
  AND2x2_ASAP7_6t_L U844 ( .A(b[11]), .B(a[12]), .Y(n579) );
  XOR2xp5r_ASAP7_6t_L U845 ( .A(n622), .B(n621), .Y(n578) );
  NOR2xp5_ASAP7_6t_L U846 ( .A(n265), .B(n516), .Y(n622) );
  AND2x2_ASAP7_6t_L U847 ( .A(a[11]), .B(b[12]), .Y(n621) );
  INVx1_ASAP7_6t_L U848 ( .A(n617), .Y(n615) );
  OAI22xp5_ASAP7_6t_L U849 ( .A1(n623), .A2(n624), .B1(n576), .B2(n577), .Y(
        n617) );
  NAND2xp5R_ASAP7_6t_L U850 ( .A(a[9]), .B(b[14]), .Y(n577) );
  XOR2xp5r_ASAP7_6t_L U851 ( .A(n625), .B(n624), .Y(n576) );
  INVx1_ASAP7_6t_L U852 ( .A(n623), .Y(n625) );
  NAND2xp5R_ASAP7_6t_L U853 ( .A(a[8]), .B(b[15]), .Y(n624) );
  AOI22xp25_ASAP7_6t_L U854 ( .A1(n626), .A2(n627), .B1(n590), .B2(n591), .Y(
        n623) );
  AND2x2_ASAP7_6t_L U855 ( .A(a[9]), .B(b[13]), .Y(n591) );
  XOR2xp5r_ASAP7_6t_L U856 ( .A(n626), .B(n627), .Y(n590) );
  NOR2xp5_ASAP7_6t_L U857 ( .A(n272), .B(n96), .Y(n627) );
  NOR2xp5_ASAP7_6t_L U858 ( .A(n402), .B(n409), .Y(n626) );
  AO21x1_ASAP7_6t_L U859 ( .A1(n628), .A2(n629), .B(n630), .Y(n1049) );
  NOR3x1f_ASAP7_6t_L U860 ( .A(n631), .B(n41), .C(n42), .Y(n630) );
  INVx1_ASAP7_6t_L U861 ( .A(n40), .Y(n631) );
  XOR2xp5r_ASAP7_6t_L U862 ( .A(n628), .B(n629), .Y(n40) );
  OAI22xp5_ASAP7_6t_L U863 ( .A1(n632), .A2(n633), .B1(n604), .B2(n603), .Y(
        n629) );
  XOR2xp5r_ASAP7_6t_L U864 ( .A(n634), .B(n635), .Y(n603) );
  XOR2xp5r_ASAP7_6t_L U865 ( .A(n636), .B(n632), .Y(n604) );
  INVx1_ASAP7_6t_L U866 ( .A(n636), .Y(n633) );
  OAI22xp5_ASAP7_6t_L U867 ( .A1(n637), .A2(n638), .B1(n639), .B2(n565), .Y(
        n636) );
  NAND2xp5R_ASAP7_6t_L U868 ( .A(b[10]), .B(a[15]), .Y(n565) );
  INVx1_ASAP7_6t_L U869 ( .A(n564), .Y(n639) );
  XOR2xp5r_ASAP7_6t_L U870 ( .A(n637), .B(n638), .Y(n564) );
  NAND2xp5R_ASAP7_6t_L U871 ( .A(b[12]), .B(a[13]), .Y(n638) );
  NAND2xp5R_ASAP7_6t_L U872 ( .A(b[11]), .B(a[14]), .Y(n637) );
  AOI22xp25_ASAP7_6t_L U873 ( .A1(n640), .A2(n641), .B1(n608), .B2(n607), .Y(
        n632) );
  XOR2xp5r_ASAP7_6t_L U874 ( .A(n641), .B(n640), .Y(n607) );
  XOR2xp5r_ASAP7_6t_L U875 ( .A(n642), .B(n643), .Y(n608) );
  OAI22xp5_ASAP7_6t_L U876 ( .A1(n644), .A2(n645), .B1(n611), .B2(n612), .Y(
        n641) );
  NAND2xp5R_ASAP7_6t_L U877 ( .A(b[10]), .B(a[14]), .Y(n612) );
  INVx1_ASAP7_6t_L U878 ( .A(n646), .Y(n611) );
  XOR2xp5r_ASAP7_6t_L U879 ( .A(n644), .B(n645), .Y(n646) );
  NAND2xp5R_ASAP7_6t_L U880 ( .A(b[12]), .B(a[12]), .Y(n645) );
  NAND2xp5R_ASAP7_6t_L U881 ( .A(b[11]), .B(a[13]), .Y(n644) );
  OAI22xp5_ASAP7_6t_L U882 ( .A1(n647), .A2(n648), .B1(n613), .B2(n614), .Y(
        n640) );
  NAND2xp5R_ASAP7_6t_L U883 ( .A(a[11]), .B(b[13]), .Y(n614) );
  XOR2xp5r_ASAP7_6t_L U884 ( .A(n649), .B(n648), .Y(n613) );
  NAND2xp5R_ASAP7_6t_L U885 ( .A(a[9]), .B(b[15]), .Y(n648) );
  INVx1_ASAP7_6t_L U886 ( .A(n649), .Y(n647) );
  NOR2xp5_ASAP7_6t_L U887 ( .A(n265), .B(n409), .Y(n649) );
  XOR2xp5r_ASAP7_6t_L U888 ( .A(n650), .B(n651), .Y(n628) );
  AO21x1_ASAP7_6t_L U889 ( .A1(n652), .A2(n653), .B(n654), .Y(n1050) );
  NOR3x1f_ASAP7_6t_L U890 ( .A(n516), .B(n38), .C(n41), .Y(n654) );
  XOR2xp5r_ASAP7_6t_L U891 ( .A(n652), .B(n655), .Y(n38) );
  INVx1_ASAP7_6t_L U892 ( .A(n655), .Y(n653) );
  AOI22xp25_ASAP7_6t_L U893 ( .A1(n656), .A2(n657), .B1(n650), .B2(n651), .Y(
        n655) );
  XOR2xp5r_ASAP7_6t_L U894 ( .A(n657), .B(n656), .Y(n651) );
  XOR2xp5r_ASAP7_6t_L U895 ( .A(n658), .B(n659), .Y(n650) );
  OAI22xp5_ASAP7_6t_L U896 ( .A1(n660), .A2(n661), .B1(n662), .B2(n602), .Y(
        n657) );
  NAND2xp5R_ASAP7_6t_L U897 ( .A(b[11]), .B(a[15]), .Y(n602) );
  INVx1_ASAP7_6t_L U898 ( .A(n601), .Y(n662) );
  XOR2xp5r_ASAP7_6t_L U899 ( .A(n661), .B(n660), .Y(n601) );
  NAND2xp5R_ASAP7_6t_L U900 ( .A(b[13]), .B(a[13]), .Y(n661) );
  NAND2xp5R_ASAP7_6t_L U901 ( .A(b[12]), .B(a[14]), .Y(n660) );
  OAI22xp5_ASAP7_6t_L U902 ( .A1(n663), .A2(n664), .B1(n665), .B2(n635), .Y(
        n656) );
  NAND2xp5R_ASAP7_6t_L U903 ( .A(a[12]), .B(b[14]), .Y(n635) );
  INVx1_ASAP7_6t_L U904 ( .A(n634), .Y(n665) );
  XOR2xp5r_ASAP7_6t_L U905 ( .A(n663), .B(n664), .Y(n634) );
  NAND2xp5R_ASAP7_6t_L U906 ( .A(a[11]), .B(b[15]), .Y(n664) );
  OA22x1_ASAP7_6t_L U907 ( .A1(n666), .A2(n667), .B1(n642), .B2(n643), .Y(n663) );
  NAND2xp5R_ASAP7_6t_L U908 ( .A(a[12]), .B(b[13]), .Y(n643) );
  INVx1_ASAP7_6t_L U909 ( .A(n668), .Y(n642) );
  XOR2xp5r_ASAP7_6t_L U910 ( .A(n666), .B(n667), .Y(n668) );
  NAND2xp5R_ASAP7_6t_L U911 ( .A(a[10]), .B(b[15]), .Y(n667) );
  NAND2xp5R_ASAP7_6t_L U912 ( .A(a[11]), .B(b[14]), .Y(n666) );
  XOR2xp5r_ASAP7_6t_L U913 ( .A(n669), .B(n670), .Y(n652) );
  OR2x2_ASAP7_6t_L U914 ( .A(n671), .B(n672), .Y(n1051) );
  NOR3x1f_ASAP7_6t_L U915 ( .A(n96), .B(n673), .C(n491), .Y(n672) );
  NOR3x1f_ASAP7_6t_L U916 ( .A(n36), .B(n41), .C(n409), .Y(n671) );
  INVx1_ASAP7_6t_L U917 ( .A(a[15]), .Y(n41) );
  XOR2xp5r_ASAP7_6t_L U918 ( .A(n674), .B(n673), .Y(n36) );
  OA22x1_ASAP7_6t_L U919 ( .A1(n675), .A2(n676), .B1(n669), .B2(n670), .Y(n673) );
  NAND2xp5R_ASAP7_6t_L U920 ( .A(a[14]), .B(b[14]), .Y(n670) );
  XOR2xp5r_ASAP7_6t_L U921 ( .A(n677), .B(n676), .Y(n669) );
  NAND2xp5R_ASAP7_6t_L U922 ( .A(b[15]), .B(a[13]), .Y(n676) );
  INVx1_ASAP7_6t_L U923 ( .A(n677), .Y(n675) );
  OAI22xp5_ASAP7_6t_L U924 ( .A1(n678), .A2(n679), .B1(n658), .B2(n659), .Y(
        n677) );
  NAND2xp5R_ASAP7_6t_L U925 ( .A(b[13]), .B(a[14]), .Y(n659) );
  XOR2xp5r_ASAP7_6t_L U926 ( .A(n680), .B(n679), .Y(n658) );
  INVx1_ASAP7_6t_L U927 ( .A(n678), .Y(n680) );
  NAND2xp5R_ASAP7_6t_L U928 ( .A(a[12]), .B(b[15]), .Y(n679) );
  NAND2xp5R_ASAP7_6t_L U929 ( .A(a[13]), .B(b[14]), .Y(n678) );
  NOR2xp5_ASAP7_6t_L U930 ( .A(n491), .B(n96), .Y(n674) );
  INVx1_ASAP7_6t_L U931 ( .A(b[15]), .Y(n96) );
  INVx1_ASAP7_6t_L U932 ( .A(n1119), .Y(n1052) );
  INVx1_ASAP7_6t_L U933 ( .A(n1118), .Y(out[14]) );
  OAI22xp5_ASAP7_6t_L U934 ( .A1(n681), .A2(n682), .B1(n67), .B2(n68), .Y(
        n1054) );
  XOR2xp5r_ASAP7_6t_L U935 ( .A(n683), .B(n681), .Y(n68) );
  XOR2xp5r_ASAP7_6t_L U936 ( .A(n684), .B(n159), .Y(n67) );
  XOR2xp5r_ASAP7_6t_L U937 ( .A(n162), .B(n161), .Y(n159) );
  XOR2xp5r_ASAP7_6t_L U938 ( .A(n147), .B(n148), .Y(n161) );
  XOR2xp5r_ASAP7_6t_L U939 ( .A(n149), .B(n150), .Y(n148) );
  XOR2xp5r_ASAP7_6t_L U940 ( .A(n217), .B(n216), .Y(n150) );
  XOR2xp5r_ASAP7_6t_L U941 ( .A(n220), .B(n218), .Y(n216) );
  INVx1_ASAP7_6t_L U942 ( .A(n685), .Y(n218) );
  XOR2xp5r_ASAP7_6t_L U943 ( .A(n282), .B(n283), .Y(n685) );
  NOR2xp5_ASAP7_6t_L U944 ( .A(n95), .B(n42), .Y(n283) );
  XOR2xp5r_ASAP7_6t_L U945 ( .A(n284), .B(n285), .Y(n282) );
  NOR2xp5_ASAP7_6t_L U946 ( .A(n99), .B(n516), .Y(n285) );
  INVx1_ASAP7_6t_L U947 ( .A(b[13]), .Y(n516) );
  NOR2xp5_ASAP7_6t_L U948 ( .A(n97), .B(n409), .Y(n284) );
  INVx1_ASAP7_6t_L U949 ( .A(b[14]), .Y(n409) );
  NOR3x1f_ASAP7_6t_L U950 ( .A(n686), .B(n42), .C(n99), .Y(n220) );
  XOR2xp5r_ASAP7_6t_L U951 ( .A(n687), .B(n280), .Y(n217) );
  NAND2xp5R_ASAP7_6t_L U952 ( .A(a[3]), .B(b[11]), .Y(n280) );
  NOR2xp5_ASAP7_6t_L U953 ( .A(n281), .B(n89), .Y(n687) );
  OAI22xp5_ASAP7_6t_L U954 ( .A1(n688), .A2(n689), .B1(n690), .B2(n691), .Y(
        n149) );
  INVx1_ASAP7_6t_L U955 ( .A(n692), .Y(n688) );
  XOR2xp5r_ASAP7_6t_L U956 ( .A(n212), .B(n213), .Y(n147) );
  NAND2xp5R_ASAP7_6t_L U957 ( .A(b[7]), .B(a[7]), .Y(n213) );
  XOR2xp5r_ASAP7_6t_L U958 ( .A(n693), .B(n215), .Y(n212) );
  NAND2xp5R_ASAP7_6t_L U959 ( .A(a[6]), .B(b[8]), .Y(n215) );
  INVx1_ASAP7_6t_L U960 ( .A(n214), .Y(n693) );
  NAND2xp5R_ASAP7_6t_L U961 ( .A(a[5]), .B(b[9]), .Y(n214) );
  XOR2xp5r_ASAP7_6t_L U962 ( .A(n151), .B(n152), .Y(n162) );
  XOR2xp5r_ASAP7_6t_L U963 ( .A(n694), .B(n153), .Y(n152) );
  AOI22xp25_ASAP7_6t_L U964 ( .A1(n695), .A2(n696), .B1(n697), .B2(n698), .Y(
        n153) );
  INVx1_ASAP7_6t_L U965 ( .A(n154), .Y(n694) );
  AOI22xp25_ASAP7_6t_L U966 ( .A1(n699), .A2(n700), .B1(n701), .B2(n702), .Y(
        n154) );
  AOI22xp25_ASAP7_6t_L U967 ( .A1(n703), .A2(n704), .B1(n705), .B2(n706), .Y(
        n151) );
  INVx1_ASAP7_6t_L U968 ( .A(n160), .Y(n684) );
  XOR2xp5r_ASAP7_6t_L U969 ( .A(n155), .B(n156), .Y(n160) );
  NOR2xp5_ASAP7_6t_L U970 ( .A(n90), .B(n491), .Y(n156) );
  INVx1_ASAP7_6t_L U971 ( .A(a[14]), .Y(n491) );
  XOR2xp5r_ASAP7_6t_L U972 ( .A(n157), .B(n158), .Y(n155) );
  XOR2xp5r_ASAP7_6t_L U973 ( .A(n202), .B(n203), .Y(n158) );
  NAND2xp5R_ASAP7_6t_L U974 ( .A(b[1]), .B(a[13]), .Y(n203) );
  INVx1_ASAP7_6t_L U975 ( .A(n707), .Y(n202) );
  XOR2xp5r_ASAP7_6t_L U976 ( .A(n205), .B(n204), .Y(n707) );
  NAND2xp5R_ASAP7_6t_L U977 ( .A(b[3]), .B(a[11]), .Y(n204) );
  NAND2xp5R_ASAP7_6t_L U978 ( .A(b[2]), .B(a[12]), .Y(n205) );
  XOR2xp5r_ASAP7_6t_L U979 ( .A(n208), .B(n209), .Y(n157) );
  NAND2xp5R_ASAP7_6t_L U980 ( .A(b[4]), .B(a[10]), .Y(n209) );
  XOR2xp5r_ASAP7_6t_L U981 ( .A(n708), .B(n210), .Y(n208) );
  NAND2xp5R_ASAP7_6t_L U982 ( .A(b[6]), .B(a[8]), .Y(n210) );
  INVx1_ASAP7_6t_L U983 ( .A(n211), .Y(n708) );
  NAND2xp5R_ASAP7_6t_L U984 ( .A(b[5]), .B(a[9]), .Y(n211) );
  INVx1_ASAP7_6t_L U985 ( .A(n683), .Y(n682) );
  XOR2xp5r_ASAP7_6t_L U986 ( .A(n108), .B(n109), .Y(n683) );
  XOR2xp5r_ASAP7_6t_L U987 ( .A(n164), .B(n163), .Y(n109) );
  OAI22xp5_ASAP7_6t_L U988 ( .A1(n709), .A2(n710), .B1(n711), .B2(n712), .Y(
        n163) );
  INVx1_ASAP7_6t_L U989 ( .A(n713), .Y(n711) );
  XOR2xp5r_ASAP7_6t_L U990 ( .A(n165), .B(n166), .Y(n164) );
  AO22x1_ASAP7_6t_L U991 ( .A1(n714), .A2(n715), .B1(n716), .B2(n717), .Y(n166) );
  OAI22xp5_ASAP7_6t_L U992 ( .A1(n718), .A2(n719), .B1(n720), .B2(n721), .Y(
        n165) );
  INVx1_ASAP7_6t_L U993 ( .A(n722), .Y(n721) );
  XOR2xp5r_ASAP7_6t_L U994 ( .A(n110), .B(n111), .Y(n108) );
  AO22x1_ASAP7_6t_L U995 ( .A1(n723), .A2(n724), .B1(n725), .B2(n726), .Y(n111) );
  OAI22xp5_ASAP7_6t_L U996 ( .A1(n727), .A2(n728), .B1(n729), .B2(n730), .Y(
        n110) );
  INVx1_ASAP7_6t_L U997 ( .A(n731), .Y(n728) );
  OA22x1_ASAP7_6t_L U998 ( .A1(n732), .A2(n733), .B1(n734), .B2(n735), .Y(n681) );
  INVx1_ASAP7_6t_L U999 ( .A(n736), .Y(n732) );
  INVx1_ASAP7_6t_L U1000 ( .A(n1117), .Y(n1055) );
  INVx1_ASAP7_6t_L U1001 ( .A(n1116), .Y(out[13]) );
  OAI22xp5_ASAP7_6t_L U1002 ( .A1(n737), .A2(n738), .B1(n70), .B2(n69), .Y(
        n1057) );
  INVx1_ASAP7_6t_L U1003 ( .A(n739), .Y(n69) );
  XOR2xp5r_ASAP7_6t_L U1004 ( .A(n723), .B(n724), .Y(n739) );
  XOR2xp5r_ASAP7_6t_L U1005 ( .A(n726), .B(n725), .Y(n724) );
  XOR2xp5r_ASAP7_6t_L U1006 ( .A(n715), .B(n714), .Y(n725) );
  XOR2xp5r_ASAP7_6t_L U1007 ( .A(n717), .B(n716), .Y(n714) );
  XOR2xp5r_ASAP7_6t_L U1008 ( .A(n696), .B(n695), .Y(n716) );
  XOR2xp5r_ASAP7_6t_L U1009 ( .A(n697), .B(n698), .Y(n695) );
  AND2x2_ASAP7_6t_L U1010 ( .A(a[2]), .B(b[11]), .Y(n698) );
  XOR2xp5r_ASAP7_6t_L U1011 ( .A(n686), .B(n740), .Y(n697) );
  NAND2xp5R_ASAP7_6t_L U1012 ( .A(a[1]), .B(b[12]), .Y(n740) );
  NAND2xp5R_ASAP7_6t_L U1013 ( .A(a[0]), .B(b[13]), .Y(n686) );
  NOR2xp5_ASAP7_6t_L U1014 ( .A(n345), .B(n281), .Y(n696) );
  NOR3x1f_ASAP7_6t_L U1015 ( .A(n741), .B(n265), .C(n742), .Y(n717) );
  XOR2xp5r_ASAP7_6t_L U1016 ( .A(n699), .B(n700), .Y(n715) );
  AND2x2_ASAP7_6t_L U1017 ( .A(a[6]), .B(b[7]), .Y(n700) );
  XOR2xp5r_ASAP7_6t_L U1018 ( .A(n702), .B(n701), .Y(n699) );
  AND2x2_ASAP7_6t_L U1019 ( .A(a[4]), .B(b[9]), .Y(n701) );
  NOR2xp5_ASAP7_6t_L U1020 ( .A(n344), .B(n271), .Y(n702) );
  XOR2xp5r_ASAP7_6t_L U1021 ( .A(n719), .B(n718), .Y(n726) );
  OA22x1_ASAP7_6t_L U1022 ( .A1(n743), .A2(n744), .B1(n745), .B2(n746), .Y(
        n718) );
  XOR2xp5r_ASAP7_6t_L U1023 ( .A(n720), .B(n722), .Y(n719) );
  OAI22xp5_ASAP7_6t_L U1024 ( .A1(n747), .A2(n748), .B1(n749), .B2(n750), .Y(
        n722) );
  AOI22xp25_ASAP7_6t_L U1025 ( .A1(n751), .A2(n752), .B1(n753), .B2(n754), .Y(
        n720) );
  XOR2xp5r_ASAP7_6t_L U1026 ( .A(n709), .B(n710), .Y(n723) );
  NAND2xp5R_ASAP7_6t_L U1027 ( .A(b[0]), .B(a[13]), .Y(n710) );
  XOR2xp5r_ASAP7_6t_L U1028 ( .A(n713), .B(n712), .Y(n709) );
  XOR2xp5r_ASAP7_6t_L U1029 ( .A(n692), .B(n689), .Y(n712) );
  NAND2xp5R_ASAP7_6t_L U1030 ( .A(b[1]), .B(a[12]), .Y(n689) );
  XOR2xp5r_ASAP7_6t_L U1031 ( .A(n691), .B(n690), .Y(n692) );
  NAND2xp5R_ASAP7_6t_L U1032 ( .A(b[3]), .B(a[10]), .Y(n690) );
  NAND2xp5R_ASAP7_6t_L U1033 ( .A(b[2]), .B(a[11]), .Y(n691) );
  XOR2xp5r_ASAP7_6t_L U1034 ( .A(n703), .B(n704), .Y(n713) );
  AND2x2_ASAP7_6t_L U1035 ( .A(b[4]), .B(a[9]), .Y(n704) );
  XOR2xp5r_ASAP7_6t_L U1036 ( .A(n706), .B(n705), .Y(n703) );
  NOR2xp5_ASAP7_6t_L U1037 ( .A(n331), .B(n272), .Y(n705) );
  NOR2xp5_ASAP7_6t_L U1038 ( .A(n264), .B(n402), .Y(n706) );
  XOR2xp5r_ASAP7_6t_L U1039 ( .A(n738), .B(n755), .Y(n70) );
  XOR2xp5r_ASAP7_6t_L U1040 ( .A(n736), .B(n733), .Y(n738) );
  XOR2xp5r_ASAP7_6t_L U1041 ( .A(n727), .B(n731), .Y(n733) );
  XOR2xp5r_ASAP7_6t_L U1042 ( .A(n730), .B(n729), .Y(n731) );
  AOI22xp25_ASAP7_6t_L U1043 ( .A1(n756), .A2(n757), .B1(n758), .B2(n759), .Y(
        n729) );
  AOI22xp25_ASAP7_6t_L U1044 ( .A1(n760), .A2(n761), .B1(n762), .B2(n763), .Y(
        n730) );
  OA22x1_ASAP7_6t_L U1045 ( .A1(n764), .A2(n765), .B1(n766), .B2(n767), .Y(
        n727) );
  INVx1_ASAP7_6t_L U1046 ( .A(n768), .Y(n764) );
  XOR2xp5r_ASAP7_6t_L U1047 ( .A(n734), .B(n735), .Y(n736) );
  AOI22xp25_ASAP7_6t_L U1048 ( .A1(n769), .A2(n770), .B1(n771), .B2(n772), .Y(
        n735) );
  INVx1_ASAP7_6t_L U1049 ( .A(n773), .Y(n770) );
  AOI22xp25_ASAP7_6t_L U1050 ( .A1(n774), .A2(n775), .B1(n776), .B2(n777), .Y(
        n734) );
  INVx1_ASAP7_6t_L U1051 ( .A(n755), .Y(n737) );
  OAI22xp5_ASAP7_6t_L U1052 ( .A1(n778), .A2(n779), .B1(n780), .B2(n781), .Y(
        n755) );
  INVx1_ASAP7_6t_L U1053 ( .A(n782), .Y(n778) );
  INVx1_ASAP7_6t_L U1054 ( .A(n1115), .Y(n1058) );
  INVx1_ASAP7_6t_L U1055 ( .A(n1114), .Y(out[12]) );
  OAI22xp5_ASAP7_6t_L U1056 ( .A1(n783), .A2(n784), .B1(n71), .B2(n72), .Y(
        n1060) );
  XOR2xp5r_ASAP7_6t_L U1057 ( .A(n785), .B(n784), .Y(n72) );
  XOR2xp5r_ASAP7_6t_L U1058 ( .A(n773), .B(n769), .Y(n71) );
  XOR2xp5r_ASAP7_6t_L U1059 ( .A(n772), .B(n771), .Y(n769) );
  XOR2xp5r_ASAP7_6t_L U1060 ( .A(n756), .B(n757), .Y(n771) );
  NOR3x1f_ASAP7_6t_L U1061 ( .A(n786), .B(n272), .C(n787), .Y(n757) );
  XOR2xp5r_ASAP7_6t_L U1062 ( .A(n759), .B(n758), .Y(n756) );
  OAI22xp5_ASAP7_6t_L U1063 ( .A1(n788), .A2(n789), .B1(n790), .B2(n791), .Y(
        n758) );
  INVx1_ASAP7_6t_L U1064 ( .A(n792), .Y(n788) );
  AO22x1_ASAP7_6t_L U1065 ( .A1(n793), .A2(n794), .B1(n795), .B2(n796), .Y(
        n759) );
  XOR2xp5r_ASAP7_6t_L U1066 ( .A(n760), .B(n761), .Y(n772) );
  XOR2xp5r_ASAP7_6t_L U1067 ( .A(n743), .B(n744), .Y(n761) );
  NAND2xp5R_ASAP7_6t_L U1068 ( .A(b[4]), .B(a[8]), .Y(n744) );
  INVx1_ASAP7_6t_L U1069 ( .A(n797), .Y(n743) );
  XOR2xp5r_ASAP7_6t_L U1070 ( .A(n745), .B(n746), .Y(n797) );
  NAND2xp5R_ASAP7_6t_L U1071 ( .A(b[5]), .B(a[7]), .Y(n746) );
  NAND2xp5R_ASAP7_6t_L U1072 ( .A(b[6]), .B(a[6]), .Y(n745) );
  XOR2xp5r_ASAP7_6t_L U1073 ( .A(n762), .B(n763), .Y(n760) );
  XOR2xp5r_ASAP7_6t_L U1074 ( .A(n747), .B(n748), .Y(n763) );
  NAND2xp5R_ASAP7_6t_L U1075 ( .A(a[5]), .B(b[7]), .Y(n748) );
  INVx1_ASAP7_6t_L U1076 ( .A(n798), .Y(n747) );
  XOR2xp5r_ASAP7_6t_L U1077 ( .A(n749), .B(n750), .Y(n798) );
  NAND2xp5R_ASAP7_6t_L U1078 ( .A(a[4]), .B(b[8]), .Y(n750) );
  NAND2xp5R_ASAP7_6t_L U1079 ( .A(a[3]), .B(b[9]), .Y(n749) );
  XOR2xp5r_ASAP7_6t_L U1080 ( .A(n751), .B(n752), .Y(n762) );
  NOR2xp5_ASAP7_6t_L U1081 ( .A(n95), .B(n281), .Y(n752) );
  XOR2xp5r_ASAP7_6t_L U1082 ( .A(n753), .B(n754), .Y(n751) );
  AND2x2_ASAP7_6t_L U1083 ( .A(a[1]), .B(b[11]), .Y(n754) );
  NOR2xp5_ASAP7_6t_L U1084 ( .A(n97), .B(n42), .Y(n753) );
  INVx1_ASAP7_6t_L U1085 ( .A(b[12]), .Y(n42) );
  XOR2xp5r_ASAP7_6t_L U1086 ( .A(n765), .B(n768), .Y(n773) );
  XOR2xp5r_ASAP7_6t_L U1087 ( .A(n766), .B(n767), .Y(n768) );
  NAND2xp5R_ASAP7_6t_L U1088 ( .A(b[1]), .B(a[11]), .Y(n767) );
  XOR2xp5r_ASAP7_6t_L U1089 ( .A(n799), .B(n741), .Y(n766) );
  NAND2xp5R_ASAP7_6t_L U1090 ( .A(b[3]), .B(a[9]), .Y(n741) );
  NOR2xp5_ASAP7_6t_L U1091 ( .A(n265), .B(n742), .Y(n799) );
  NAND2xp5R_ASAP7_6t_L U1092 ( .A(b[0]), .B(a[12]), .Y(n765) );
  XOR2xp5r_ASAP7_6t_L U1093 ( .A(n779), .B(n782), .Y(n784) );
  XOR2xp5r_ASAP7_6t_L U1094 ( .A(n780), .B(n781), .Y(n782) );
  AOI22xp25_ASAP7_6t_L U1095 ( .A1(n800), .A2(n801), .B1(n802), .B2(n803), .Y(
        n781) );
  AOI22xp25_ASAP7_6t_L U1096 ( .A1(n804), .A2(n805), .B1(n806), .B2(n807), .Y(
        n780) );
  INVx1_ASAP7_6t_L U1097 ( .A(n808), .Y(n804) );
  INVx1_ASAP7_6t_L U1098 ( .A(n809), .Y(n779) );
  XOR2xp5r_ASAP7_6t_L U1099 ( .A(n774), .B(n775), .Y(n809) );
  XOR2xp5r_ASAP7_6t_L U1100 ( .A(n777), .B(n776), .Y(n775) );
  OAI22xp5_ASAP7_6t_L U1101 ( .A1(n810), .A2(n811), .B1(n812), .B2(n813), .Y(
        n776) );
  INVx1_ASAP7_6t_L U1102 ( .A(n814), .Y(n813) );
  AO22x1_ASAP7_6t_L U1103 ( .A1(n815), .A2(n816), .B1(n817), .B2(n818), .Y(
        n777) );
  OAI22xp5_ASAP7_6t_L U1104 ( .A1(n819), .A2(n820), .B1(n821), .B2(n822), .Y(
        n774) );
  INVx1_ASAP7_6t_L U1105 ( .A(n785), .Y(n783) );
  OAI22xp5_ASAP7_6t_L U1106 ( .A1(n823), .A2(n824), .B1(n825), .B2(n826), .Y(
        n785) );
  INVx1_ASAP7_6t_L U1107 ( .A(n827), .Y(n825) );
  INVx1_ASAP7_6t_L U1108 ( .A(n1113), .Y(n1061) );
  INVx1_ASAP7_6t_L U1109 ( .A(n1112), .Y(out[11]) );
  OAI22xp5_ASAP7_6t_L U1110 ( .A1(n828), .A2(n829), .B1(n74), .B2(n73), .Y(
        n1063) );
  INVx1_ASAP7_6t_L U1111 ( .A(n830), .Y(n73) );
  XOR2xp5r_ASAP7_6t_L U1112 ( .A(n800), .B(n801), .Y(n830) );
  XOR2xp5r_ASAP7_6t_L U1113 ( .A(n802), .B(n803), .Y(n801) );
  XOR2xp5r_ASAP7_6t_L U1114 ( .A(n811), .B(n810), .Y(n803) );
  XOR2xp5r_ASAP7_6t_L U1115 ( .A(n792), .B(n789), .Y(n810) );
  NAND2xp5R_ASAP7_6t_L U1116 ( .A(a[2]), .B(b[9]), .Y(n789) );
  XOR2xp5r_ASAP7_6t_L U1117 ( .A(n790), .B(n791), .Y(n792) );
  NAND2xp5R_ASAP7_6t_L U1118 ( .A(a[1]), .B(b[10]), .Y(n791) );
  NAND2xp5R_ASAP7_6t_L U1119 ( .A(a[0]), .B(b[11]), .Y(n790) );
  XOR2xp5r_ASAP7_6t_L U1120 ( .A(n812), .B(n814), .Y(n811) );
  NOR3x1f_ASAP7_6t_L U1121 ( .A(n831), .B(n331), .C(n89), .Y(n814) );
  AOI22xp25_ASAP7_6t_L U1122 ( .A1(n832), .A2(n833), .B1(n834), .B2(n835), .Y(
        n812) );
  XOR2xp5r_ASAP7_6t_L U1123 ( .A(n816), .B(n815), .Y(n802) );
  XOR2xp5r_ASAP7_6t_L U1124 ( .A(n818), .B(n817), .Y(n815) );
  XOR2xp5r_ASAP7_6t_L U1125 ( .A(n793), .B(n794), .Y(n817) );
  NOR2xp5_ASAP7_6t_L U1126 ( .A(n344), .B(n331), .Y(n794) );
  XOR2xp5r_ASAP7_6t_L U1127 ( .A(n795), .B(n796), .Y(n793) );
  AND2x2_ASAP7_6t_L U1128 ( .A(a[4]), .B(b[7]), .Y(n796) );
  NOR2xp5_ASAP7_6t_L U1129 ( .A(n345), .B(n271), .Y(n795) );
  XOR2xp5r_ASAP7_6t_L U1130 ( .A(n836), .B(n786), .Y(n818) );
  NAND2xp5R_ASAP7_6t_L U1131 ( .A(b[5]), .B(a[6]), .Y(n786) );
  NAND2xp5R_ASAP7_6t_L U1132 ( .A(a[7]), .B(b[4]), .Y(n836) );
  NOR2xp5_ASAP7_6t_L U1133 ( .A(n837), .B(n402), .Y(n816) );
  XOR2xp5r_ASAP7_6t_L U1134 ( .A(n819), .B(n820), .Y(n800) );
  NAND2xp5R_ASAP7_6t_L U1135 ( .A(b[0]), .B(a[11]), .Y(n820) );
  XOR2xp5r_ASAP7_6t_L U1136 ( .A(n838), .B(n822), .Y(n819) );
  NAND2xp5R_ASAP7_6t_L U1137 ( .A(b[1]), .B(a[10]), .Y(n822) );
  INVx1_ASAP7_6t_L U1138 ( .A(n821), .Y(n838) );
  NAND2xp5R_ASAP7_6t_L U1139 ( .A(b[2]), .B(a[9]), .Y(n821) );
  XOR2xp5r_ASAP7_6t_L U1140 ( .A(n828), .B(n839), .Y(n74) );
  INVx1_ASAP7_6t_L U1141 ( .A(n839), .Y(n829) );
  XOR2xp5r_ASAP7_6t_L U1142 ( .A(n824), .B(n823), .Y(n839) );
  XOR2xp5r_ASAP7_6t_L U1143 ( .A(n827), .B(n826), .Y(n823) );
  AOI22xp25_ASAP7_6t_L U1144 ( .A1(n840), .A2(n841), .B1(n842), .B2(n843), .Y(
        n826) );
  OAI22xp5_ASAP7_6t_L U1145 ( .A1(n844), .A2(n845), .B1(n846), .B2(n847), .Y(
        n827) );
  XOR2xp5r_ASAP7_6t_L U1146 ( .A(n808), .B(n805), .Y(n824) );
  XOR2xp5r_ASAP7_6t_L U1147 ( .A(n807), .B(n806), .Y(n805) );
  OAI22xp5_ASAP7_6t_L U1148 ( .A1(n848), .A2(n849), .B1(n850), .B2(n851), .Y(
        n806) );
  INVx1_ASAP7_6t_L U1149 ( .A(n852), .Y(n851) );
  OAI22xp5_ASAP7_6t_L U1150 ( .A1(n853), .A2(n854), .B1(n855), .B2(n856), .Y(
        n807) );
  AOI22xp25_ASAP7_6t_L U1151 ( .A1(n857), .A2(n858), .B1(n859), .B2(n860), .Y(
        n808) );
  AOI22xp25_ASAP7_6t_L U1152 ( .A1(n861), .A2(n862), .B1(n863), .B2(n864), .Y(
        n828) );
  INVx1_ASAP7_6t_L U1153 ( .A(n1111), .Y(n1064) );
  INVx1_ASAP7_6t_L U1154 ( .A(n1110), .Y(out[10]) );
  OAI22xp5_ASAP7_6t_L U1155 ( .A1(n865), .A2(n866), .B1(n75), .B2(n76), .Y(
        n1066) );
  XOR2xp5r_ASAP7_6t_L U1156 ( .A(n867), .B(n865), .Y(n76) );
  XOR2xp5r_ASAP7_6t_L U1157 ( .A(n868), .B(n840), .Y(n75) );
  XOR2xp5r_ASAP7_6t_L U1158 ( .A(n843), .B(n842), .Y(n840) );
  XOR2xp5r_ASAP7_6t_L U1159 ( .A(n849), .B(n848), .Y(n842) );
  XOR2xp5r_ASAP7_6t_L U1160 ( .A(n852), .B(n850), .Y(n848) );
  INVx1_ASAP7_6t_L U1161 ( .A(n869), .Y(n850) );
  XOR2xp5r_ASAP7_6t_L U1162 ( .A(n832), .B(n833), .Y(n869) );
  NOR2xp5_ASAP7_6t_L U1163 ( .A(n95), .B(n271), .Y(n833) );
  XOR2xp5r_ASAP7_6t_L U1164 ( .A(n834), .B(n835), .Y(n832) );
  AND2x2_ASAP7_6t_L U1165 ( .A(a[1]), .B(b[9]), .Y(n835) );
  NOR2xp5_ASAP7_6t_L U1166 ( .A(n97), .B(n281), .Y(n834) );
  INVx1_ASAP7_6t_L U1167 ( .A(b[10]), .Y(n281) );
  NOR3x1f_ASAP7_6t_L U1168 ( .A(n870), .B(n271), .C(n99), .Y(n852) );
  XOR2xp5r_ASAP7_6t_L U1169 ( .A(n871), .B(n831), .Y(n849) );
  NAND2xp5R_ASAP7_6t_L U1170 ( .A(a[3]), .B(b[7]), .Y(n831) );
  NOR2xp5_ASAP7_6t_L U1171 ( .A(n331), .B(n89), .Y(n871) );
  XOR2xp5r_ASAP7_6t_L U1172 ( .A(n853), .B(n854), .Y(n843) );
  NAND2xp5R_ASAP7_6t_L U1173 ( .A(b[3]), .B(a[7]), .Y(n854) );
  XOR2xp5r_ASAP7_6t_L U1174 ( .A(n872), .B(n855), .Y(n853) );
  NAND2xp5R_ASAP7_6t_L U1175 ( .A(b[5]), .B(a[5]), .Y(n855) );
  INVx1_ASAP7_6t_L U1176 ( .A(n856), .Y(n872) );
  NAND2xp5R_ASAP7_6t_L U1177 ( .A(b[4]), .B(a[6]), .Y(n856) );
  INVx1_ASAP7_6t_L U1178 ( .A(n841), .Y(n868) );
  XOR2xp5r_ASAP7_6t_L U1179 ( .A(n857), .B(n858), .Y(n841) );
  NOR2xp5_ASAP7_6t_L U1180 ( .A(n90), .B(n265), .Y(n858) );
  INVx1_ASAP7_6t_L U1181 ( .A(a[10]), .Y(n265) );
  XOR2xp5r_ASAP7_6t_L U1182 ( .A(n859), .B(n860), .Y(n857) );
  AND2x2_ASAP7_6t_L U1183 ( .A(b[1]), .B(a[9]), .Y(n860) );
  NOR2xp5_ASAP7_6t_L U1184 ( .A(n742), .B(n402), .Y(n859) );
  INVx1_ASAP7_6t_L U1185 ( .A(n867), .Y(n866) );
  XOR2xp5r_ASAP7_6t_L U1186 ( .A(n861), .B(n862), .Y(n867) );
  XOR2xp5r_ASAP7_6t_L U1187 ( .A(n844), .B(n845), .Y(n862) );
  INVx1_ASAP7_6t_L U1188 ( .A(n873), .Y(n845) );
  XOR2xp5r_ASAP7_6t_L U1189 ( .A(n847), .B(n846), .Y(n873) );
  AOI22xp25_ASAP7_6t_L U1190 ( .A1(n874), .A2(n875), .B1(n876), .B2(n877), .Y(
        n846) );
  AOI22xp25_ASAP7_6t_L U1191 ( .A1(n878), .A2(n879), .B1(n880), .B2(n881), .Y(
        n847) );
  AOI22xp25_ASAP7_6t_L U1192 ( .A1(n882), .A2(n883), .B1(n884), .B2(n885), .Y(
        n844) );
  XOR2xp5r_ASAP7_6t_L U1193 ( .A(n863), .B(n864), .Y(n861) );
  AO22x1_ASAP7_6t_L U1194 ( .A1(n886), .A2(n887), .B1(n888), .B2(n889), .Y(
        n864) );
  AO22x1_ASAP7_6t_L U1195 ( .A1(n890), .A2(n891), .B1(n892), .B2(n893), .Y(
        n863) );
  AOI22xp25_ASAP7_6t_L U1196 ( .A1(n894), .A2(n895), .B1(n896), .B2(n897), .Y(
        n865) );
  INVx1_ASAP7_6t_L U1197 ( .A(n1109), .Y(n1067) );
  INVx1_ASAP7_6t_L U1198 ( .A(n1108), .Y(out[9]) );
  OAI22xp5_ASAP7_6t_L U1199 ( .A1(n898), .A2(n899), .B1(n77), .B2(n78), .Y(
        n1069) );
  XOR2xp5r_ASAP7_6t_L U1200 ( .A(n898), .B(n900), .Y(n78) );
  XOR2xp5r_ASAP7_6t_L U1201 ( .A(n901), .B(n886), .Y(n77) );
  XOR2xp5r_ASAP7_6t_L U1202 ( .A(n889), .B(n888), .Y(n886) );
  XOR2xp5r_ASAP7_6t_L U1203 ( .A(n875), .B(n874), .Y(n888) );
  XOR2xp5r_ASAP7_6t_L U1204 ( .A(n876), .B(n877), .Y(n874) );
  AND2x2_ASAP7_6t_L U1205 ( .A(a[2]), .B(b[7]), .Y(n877) );
  XOR2xp5r_ASAP7_6t_L U1206 ( .A(n870), .B(n902), .Y(n876) );
  NAND2xp5R_ASAP7_6t_L U1207 ( .A(a[1]), .B(b[8]), .Y(n902) );
  NAND2xp5R_ASAP7_6t_L U1208 ( .A(a[0]), .B(b[9]), .Y(n870) );
  NOR2xp5_ASAP7_6t_L U1209 ( .A(n345), .B(n331), .Y(n875) );
  XOR2xp5r_ASAP7_6t_L U1210 ( .A(n878), .B(n879), .Y(n889) );
  AND2x2_ASAP7_6t_L U1211 ( .A(b[3]), .B(a[6]), .Y(n879) );
  XOR2xp5r_ASAP7_6t_L U1212 ( .A(n881), .B(n880), .Y(n878) );
  NOR2xp5_ASAP7_6t_L U1213 ( .A(n89), .B(n264), .Y(n880) );
  NOR2xp5_ASAP7_6t_L U1214 ( .A(n787), .B(n344), .Y(n881) );
  INVx1_ASAP7_6t_L U1215 ( .A(n887), .Y(n901) );
  XOR2xp5r_ASAP7_6t_L U1216 ( .A(n882), .B(n883), .Y(n887) );
  AND2x2_ASAP7_6t_L U1217 ( .A(b[0]), .B(a[9]), .Y(n883) );
  XOR2xp5r_ASAP7_6t_L U1218 ( .A(n884), .B(n885), .Y(n882) );
  NOR2xp5_ASAP7_6t_L U1219 ( .A(n98), .B(n402), .Y(n885) );
  INVx1_ASAP7_6t_L U1220 ( .A(a[8]), .Y(n402) );
  NOR2xp5_ASAP7_6t_L U1221 ( .A(n742), .B(n272), .Y(n884) );
  INVx1_ASAP7_6t_L U1222 ( .A(n900), .Y(n899) );
  XOR2xp5r_ASAP7_6t_L U1223 ( .A(n895), .B(n894), .Y(n900) );
  XOR2xp5r_ASAP7_6t_L U1224 ( .A(n897), .B(n896), .Y(n894) );
  OAI22xp5_ASAP7_6t_L U1225 ( .A1(n903), .A2(n904), .B1(n905), .B2(n906), .Y(
        n896) );
  INVx1_ASAP7_6t_L U1226 ( .A(n907), .Y(n905) );
  AO22x1_ASAP7_6t_L U1227 ( .A1(n908), .A2(n909), .B1(n910), .B2(n911), .Y(
        n897) );
  INVx1_ASAP7_6t_L U1228 ( .A(n912), .Y(n909) );
  XOR2xp5r_ASAP7_6t_L U1229 ( .A(n890), .B(n891), .Y(n895) );
  NOR3x1f_ASAP7_6t_L U1230 ( .A(n913), .B(n272), .C(n98), .Y(n891) );
  XOR2xp5r_ASAP7_6t_L U1231 ( .A(n892), .B(n893), .Y(n890) );
  OAI22xp5_ASAP7_6t_L U1232 ( .A1(n914), .A2(n915), .B1(n916), .B2(n917), .Y(
        n893) );
  AO22x1_ASAP7_6t_L U1233 ( .A1(n918), .A2(n919), .B1(n920), .B2(n921), .Y(
        n892) );
  AOI22xp25_ASAP7_6t_L U1234 ( .A1(n922), .A2(n923), .B1(n924), .B2(n925), .Y(
        n898) );
  INVx1_ASAP7_6t_L U1235 ( .A(n1107), .Y(n1070) );
  INVx1_ASAP7_6t_L U1236 ( .A(n1106), .Y(out[8]) );
  OAI22xp5_ASAP7_6t_L U1237 ( .A1(n926), .A2(n927), .B1(n79), .B2(n80), .Y(
        n1072) );
  XOR2xp5r_ASAP7_6t_L U1238 ( .A(n926), .B(n928), .Y(n80) );
  XOR2xp5r_ASAP7_6t_L U1239 ( .A(n912), .B(n908), .Y(n79) );
  XOR2xp5r_ASAP7_6t_L U1240 ( .A(n911), .B(n910), .Y(n908) );
  XOR2xp5r_ASAP7_6t_L U1241 ( .A(n914), .B(n915), .Y(n910) );
  NAND2xp5R_ASAP7_6t_L U1242 ( .A(b[3]), .B(a[5]), .Y(n915) );
  XOR2xp5r_ASAP7_6t_L U1243 ( .A(n929), .B(n917), .Y(n914) );
  NAND2xp5R_ASAP7_6t_L U1244 ( .A(b[4]), .B(a[4]), .Y(n917) );
  INVx1_ASAP7_6t_L U1245 ( .A(n916), .Y(n929) );
  NAND2xp5R_ASAP7_6t_L U1246 ( .A(a[3]), .B(b[5]), .Y(n916) );
  XOR2xp5r_ASAP7_6t_L U1247 ( .A(n930), .B(n913), .Y(n911) );
  NAND2xp5R_ASAP7_6t_L U1248 ( .A(b[2]), .B(a[6]), .Y(n913) );
  NAND2xp5R_ASAP7_6t_L U1249 ( .A(a[7]), .B(b[1]), .Y(n930) );
  NAND2xp5R_ASAP7_6t_L U1250 ( .A(b[0]), .B(a[8]), .Y(n912) );
  INVx1_ASAP7_6t_L U1251 ( .A(n928), .Y(n927) );
  XOR2xp5r_ASAP7_6t_L U1252 ( .A(n922), .B(n923), .Y(n928) );
  XOR2xp5r_ASAP7_6t_L U1253 ( .A(n904), .B(n903), .Y(n923) );
  INVx1_ASAP7_6t_L U1254 ( .A(n931), .Y(n903) );
  XOR2xp5r_ASAP7_6t_L U1255 ( .A(n918), .B(n919), .Y(n931) );
  NOR2xp5_ASAP7_6t_L U1256 ( .A(n95), .B(n331), .Y(n919) );
  INVx1_ASAP7_6t_L U1257 ( .A(b[6]), .Y(n331) );
  XOR2xp5r_ASAP7_6t_L U1258 ( .A(n920), .B(n921), .Y(n918) );
  AND2x2_ASAP7_6t_L U1259 ( .A(a[1]), .B(b[7]), .Y(n921) );
  NOR2xp5_ASAP7_6t_L U1260 ( .A(n97), .B(n271), .Y(n920) );
  INVx1_ASAP7_6t_L U1261 ( .A(b[8]), .Y(n271) );
  XOR2xp5r_ASAP7_6t_L U1262 ( .A(n907), .B(n906), .Y(n904) );
  NAND3xp33R_ASAP7_6t_L U1263 ( .A(n932), .B(a[4]), .C(b[3]), .Y(n906) );
  OAI22xp5_ASAP7_6t_L U1264 ( .A1(n933), .A2(n934), .B1(n935), .B2(n936), .Y(
        n907) );
  INVx1_ASAP7_6t_L U1265 ( .A(n937), .Y(n933) );
  XOR2xp5r_ASAP7_6t_L U1266 ( .A(n925), .B(n924), .Y(n922) );
  OAI22xp5_ASAP7_6t_L U1267 ( .A1(n938), .A2(n939), .B1(n940), .B2(n941), .Y(
        n924) );
  INVx1_ASAP7_6t_L U1268 ( .A(n942), .Y(n941) );
  AO22x1_ASAP7_6t_L U1269 ( .A1(n943), .A2(n944), .B1(n945), .B2(n946), .Y(
        n925) );
  AOI22xp25_ASAP7_6t_L U1270 ( .A1(n947), .A2(n948), .B1(n949), .B2(n950), .Y(
        n926) );
  INVx1_ASAP7_6t_L U1271 ( .A(n1105), .Y(n1073) );
  INVx1_ASAP7_6t_L U1272 ( .A(n1104), .Y(out[7]) );
  OAI22xp5_ASAP7_6t_L U1273 ( .A1(n951), .A2(n952), .B1(n81), .B2(n82), .Y(
        n1075) );
  XOR2xp5r_ASAP7_6t_L U1274 ( .A(n951), .B(n953), .Y(n82) );
  INVx1_ASAP7_6t_L U1275 ( .A(n954), .Y(n81) );
  XOR2xp5r_ASAP7_6t_L U1276 ( .A(n943), .B(n944), .Y(n954) );
  NOR2xp5_ASAP7_6t_L U1277 ( .A(n90), .B(n272), .Y(n944) );
  INVx1_ASAP7_6t_L U1278 ( .A(a[7]), .Y(n272) );
  XOR2xp5r_ASAP7_6t_L U1279 ( .A(n945), .B(n946), .Y(n943) );
  AND2x2_ASAP7_6t_L U1280 ( .A(b[1]), .B(a[6]), .Y(n946) );
  NOR2xp5_ASAP7_6t_L U1281 ( .A(n742), .B(n344), .Y(n945) );
  INVx1_ASAP7_6t_L U1282 ( .A(n953), .Y(n952) );
  XOR2xp5r_ASAP7_6t_L U1283 ( .A(n948), .B(n947), .Y(n953) );
  XOR2xp5r_ASAP7_6t_L U1284 ( .A(n950), .B(n949), .Y(n947) );
  AO22x1_ASAP7_6t_L U1285 ( .A1(n955), .A2(n956), .B1(n957), .B2(n958), .Y(
        n949) );
  AO22x1_ASAP7_6t_L U1286 ( .A1(n959), .A2(n960), .B1(n961), .B2(n962), .Y(
        n950) );
  XOR2xp5r_ASAP7_6t_L U1287 ( .A(n939), .B(n938), .Y(n948) );
  XOR2xp5r_ASAP7_6t_L U1288 ( .A(n942), .B(n940), .Y(n938) );
  XOR2xp5r_ASAP7_6t_L U1289 ( .A(n937), .B(n934), .Y(n940) );
  NAND2xp5R_ASAP7_6t_L U1290 ( .A(a[2]), .B(b[5]), .Y(n934) );
  XOR2xp5r_ASAP7_6t_L U1291 ( .A(n935), .B(n936), .Y(n937) );
  NAND2xp5R_ASAP7_6t_L U1292 ( .A(a[1]), .B(b[6]), .Y(n936) );
  NAND2xp5R_ASAP7_6t_L U1293 ( .A(a[0]), .B(b[7]), .Y(n935) );
  NOR3x1f_ASAP7_6t_L U1294 ( .A(n963), .B(n264), .C(n99), .Y(n942) );
  XOR2xp5r_ASAP7_6t_L U1295 ( .A(n932), .B(n964), .Y(n939) );
  NAND2xp5R_ASAP7_6t_L U1296 ( .A(b[3]), .B(a[4]), .Y(n964) );
  NOR2xp5_ASAP7_6t_L U1297 ( .A(n787), .B(n345), .Y(n932) );
  AOI22xp25_ASAP7_6t_L U1298 ( .A1(n965), .A2(n966), .B1(n967), .B2(n968), .Y(
        n951) );
  INVx1_ASAP7_6t_L U1299 ( .A(n1103), .Y(n1076) );
  INVx1_ASAP7_6t_L U1300 ( .A(n1102), .Y(out[6]) );
  OAI22xp5_ASAP7_6t_L U1301 ( .A1(n969), .A2(n970), .B1(n83), .B2(n84), .Y(
        n1078) );
  XOR2xp5r_ASAP7_6t_L U1302 ( .A(n969), .B(n971), .Y(n84) );
  XOR2xp5r_ASAP7_6t_L U1303 ( .A(n972), .B(n960), .Y(n83) );
  AND2x2_ASAP7_6t_L U1304 ( .A(b[0]), .B(a[6]), .Y(n960) );
  INVx1_ASAP7_6t_L U1305 ( .A(n959), .Y(n972) );
  XOR2xp5r_ASAP7_6t_L U1306 ( .A(n962), .B(n961), .Y(n959) );
  NOR2xp5_ASAP7_6t_L U1307 ( .A(n742), .B(n89), .Y(n961) );
  NOR2xp5_ASAP7_6t_L U1308 ( .A(n98), .B(n344), .Y(n962) );
  INVx1_ASAP7_6t_L U1309 ( .A(n971), .Y(n970) );
  XOR2xp5r_ASAP7_6t_L U1310 ( .A(n966), .B(n965), .Y(n971) );
  XOR2xp5r_ASAP7_6t_L U1311 ( .A(n956), .B(n955), .Y(n965) );
  XOR2xp5r_ASAP7_6t_L U1312 ( .A(n957), .B(n958), .Y(n955) );
  NOR2xp5_ASAP7_6t_L U1313 ( .A(n95), .B(n787), .Y(n958) );
  XOR2xp5r_ASAP7_6t_L U1314 ( .A(n963), .B(n973), .Y(n957) );
  NAND2xp5R_ASAP7_6t_L U1315 ( .A(a[1]), .B(b[5]), .Y(n973) );
  NAND2xp5R_ASAP7_6t_L U1316 ( .A(a[0]), .B(b[6]), .Y(n963) );
  NOR2xp5_ASAP7_6t_L U1317 ( .A(n837), .B(n345), .Y(n956) );
  XOR2xp5r_ASAP7_6t_L U1318 ( .A(n967), .B(n968), .Y(n966) );
  NOR3x1f_ASAP7_6t_L U1319 ( .A(n974), .B(n89), .C(n98), .Y(n968) );
  AO22x1_ASAP7_6t_L U1320 ( .A1(n975), .A2(n976), .B1(n977), .B2(n978), .Y(
        n967) );
  AOI22xp25_ASAP7_6t_L U1321 ( .A1(n979), .A2(n980), .B1(n981), .B2(n982), .Y(
        n969) );
  INVx1_ASAP7_6t_L U1322 ( .A(n1101), .Y(n1079) );
  INVx1_ASAP7_6t_L U1323 ( .A(n1100), .Y(out[5]) );
  AO21x1_ASAP7_6t_L U1324 ( .A1(n983), .A2(n984), .B(n985), .Y(n1081) );
  NOR3x1f_ASAP7_6t_L U1325 ( .A(n86), .B(n344), .C(n90), .Y(n985) );
  INVx1_ASAP7_6t_L U1326 ( .A(a[5]), .Y(n344) );
  XOR2xp5r_ASAP7_6t_L U1327 ( .A(n986), .B(n983), .Y(n86) );
  INVx1_ASAP7_6t_L U1328 ( .A(n986), .Y(n984) );
  AOI22xp25_ASAP7_6t_L U1329 ( .A1(n987), .A2(n988), .B1(n989), .B2(n990), .Y(
        n986) );
  XOR2xp5r_ASAP7_6t_L U1330 ( .A(n980), .B(n979), .Y(n983) );
  XOR2xp5r_ASAP7_6t_L U1331 ( .A(n982), .B(n981), .Y(n979) );
  XOR2xp5r_ASAP7_6t_L U1332 ( .A(n975), .B(n976), .Y(n981) );
  NOR2xp5_ASAP7_6t_L U1333 ( .A(n837), .B(n95), .Y(n976) );
  XOR2xp5r_ASAP7_6t_L U1334 ( .A(n977), .B(n978), .Y(n975) );
  NOR2xp5_ASAP7_6t_L U1335 ( .A(n99), .B(n787), .Y(n978) );
  INVx1_ASAP7_6t_L U1336 ( .A(b[4]), .Y(n787) );
  NOR2xp5_ASAP7_6t_L U1337 ( .A(n97), .B(n264), .Y(n977) );
  INVx1_ASAP7_6t_L U1338 ( .A(b[5]), .Y(n264) );
  INVx1_ASAP7_6t_L U1339 ( .A(a[0]), .Y(n97) );
  NOR3x1f_ASAP7_6t_L U1340 ( .A(n991), .B(n837), .C(n99), .Y(n982) );
  INVx1_ASAP7_6t_L U1341 ( .A(b[3]), .Y(n837) );
  XOR2xp5r_ASAP7_6t_L U1342 ( .A(n992), .B(n974), .Y(n980) );
  NAND2xp5R_ASAP7_6t_L U1343 ( .A(b[2]), .B(a[3]), .Y(n974) );
  NAND2xp5R_ASAP7_6t_L U1344 ( .A(a[4]), .B(b[1]), .Y(n992) );
  INVx1_ASAP7_6t_L U1345 ( .A(n1099), .Y(n1082) );
  INVx1_ASAP7_6t_L U1346 ( .A(n1098), .Y(out[4]) );
  AO21x1_ASAP7_6t_L U1347 ( .A1(n993), .A2(n994), .B(n995), .Y(n1084) );
  NOR3x1f_ASAP7_6t_L U1348 ( .A(n90), .B(n996), .C(n89), .Y(n995) );
  INVx1_ASAP7_6t_L U1349 ( .A(a[4]), .Y(n89) );
  INVx1_ASAP7_6t_L U1350 ( .A(n88), .Y(n996) );
  XOR2xp5r_ASAP7_6t_L U1351 ( .A(n993), .B(n994), .Y(n88) );
  XOR2xp5r_ASAP7_6t_L U1352 ( .A(n988), .B(n987), .Y(n994) );
  XOR2xp5r_ASAP7_6t_L U1353 ( .A(n989), .B(n990), .Y(n987) );
  NOR2xp5_ASAP7_6t_L U1354 ( .A(n742), .B(n95), .Y(n990) );
  XOR2xp5r_ASAP7_6t_L U1355 ( .A(n991), .B(n997), .Y(n989) );
  NAND2xp5R_ASAP7_6t_L U1356 ( .A(a[1]), .B(b[3]), .Y(n997) );
  NAND2xp5R_ASAP7_6t_L U1357 ( .A(a[0]), .B(b[4]), .Y(n991) );
  NOR2xp5_ASAP7_6t_L U1358 ( .A(n98), .B(n345), .Y(n988) );
  NOR3x1f_ASAP7_6t_L U1359 ( .A(n998), .B(n99), .C(n742), .Y(n993) );
  INVx1_ASAP7_6t_L U1360 ( .A(b[2]), .Y(n742) );
  INVx1_ASAP7_6t_L U1361 ( .A(n1097), .Y(n1085) );
  INVx1_ASAP7_6t_L U1362 ( .A(n1096), .Y(out[3]) );
  OR2x2_ASAP7_6t_L U1363 ( .A(n999), .B(n1000), .Y(n1087) );
  NOR3x1f_ASAP7_6t_L U1364 ( .A(n98), .B(n1001), .C(n95), .Y(n1000) );
  INVx1_ASAP7_6t_L U1365 ( .A(a[2]), .Y(n95) );
  INVx1_ASAP7_6t_L U1366 ( .A(n1002), .Y(n1001) );
  NOR3x1f_ASAP7_6t_L U1367 ( .A(n90), .B(n91), .C(n345), .Y(n999) );
  INVx1_ASAP7_6t_L U1368 ( .A(a[3]), .Y(n345) );
  XOR2xp5r_ASAP7_6t_L U1369 ( .A(n1002), .B(n1003), .Y(n91) );
  NAND2xp5R_ASAP7_6t_L U1370 ( .A(b[1]), .B(a[2]), .Y(n1003) );
  XOR2xp5r_ASAP7_6t_L U1371 ( .A(n998), .B(n1004), .Y(n1002) );
  NAND2xp5R_ASAP7_6t_L U1372 ( .A(b[2]), .B(a[1]), .Y(n1004) );
  NAND2xp5R_ASAP7_6t_L U1373 ( .A(a[0]), .B(b[3]), .Y(n998) );
  INVx1_ASAP7_6t_L U1374 ( .A(b[0]), .Y(n90) );
  INVx1_ASAP7_6t_L U1375 ( .A(n1095), .Y(n1088) );
  INVx1_ASAP7_6t_L U1376 ( .A(n1094), .Y(out[2]) );
  INVx1_ASAP7_6t_L U1377 ( .A(n1093), .Y(n1090) );
  INVx1_ASAP7_6t_L U1378 ( .A(n1092), .Y(out[1]) );
  NOR3x1f_ASAP7_6t_L U1379 ( .A(n94), .B(n99), .C(n98), .Y(c_182_) );
  INVx1_ASAP7_6t_L U1380 ( .A(b[1]), .Y(n98) );
  INVx1_ASAP7_6t_L U1381 ( .A(a[1]), .Y(n99) );
  NAND2xp5R_ASAP7_6t_L U1382 ( .A(a[0]), .B(b[2]), .Y(n94) );
endmodule

