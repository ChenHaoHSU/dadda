
module DADDA_8x8_52 ( a, b, out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] out;
  wire   n19, n20, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n239, n241, n243, n245, n247, n249, n251, n253, n254, n256,
         n258, n260, n261, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286;
  wire   [16:1] p;
  wire   [21:9] s;
  wire   [20:9] c;

  FAxp33_ASAP7_6t_L add_78_U1_1 ( .A(s[9]), .B(p[16]), .CI(n19), .CON(n264), 
        .SN(n263) );
  FAxp33_ASAP7_6t_L add_78_U1_2 ( .A(n260), .B(c[9]), .CI(n261), .CON(n266), 
        .SN(n265) );
  FAxp33_ASAP7_6t_L add_78_U1_4 ( .A(s[12]), .B(c[11]), .CI(n20), .CON(n268), 
        .SN(n267) );
  FAxp33_ASAP7_6t_L add_78_U1_5 ( .A(s[13]), .B(c[12]), .CI(n256), .CON(n270), 
        .SN(n269) );
  FAxp33_ASAP7_6t_L add_78_U1_6 ( .A(s[14]), .B(c[13]), .CI(n254), .CON(n272), 
        .SN(n271) );
  FAxp33_ASAP7_6t_L add_78_U1_7 ( .A(s[15]), .B(c[14]), .CI(n251), .CON(n274), 
        .SN(n273) );
  FAxp33_ASAP7_6t_L add_78_U1_8 ( .A(s[16]), .B(c[15]), .CI(n249), .CON(n276), 
        .SN(n275) );
  FAxp33_ASAP7_6t_L add_78_U1_9 ( .A(s[17]), .B(c[16]), .CI(n247), .CON(n278), 
        .SN(n277) );
  FAxp33_ASAP7_6t_L add_78_U1_10 ( .A(s[18]), .B(c[17]), .CI(n245), .CON(n280), 
        .SN(n279) );
  FAxp33_ASAP7_6t_L add_78_U1_11 ( .A(s[19]), .B(c[18]), .CI(n243), .CON(n282), 
        .SN(n281) );
  FAxp33_ASAP7_6t_L add_78_U1_12 ( .A(s[20]), .B(c[19]), .CI(n241), .CON(n284), 
        .SN(n283) );
  FAxp33_ASAP7_6t_L add_78_U1_13 ( .A(s[21]), .B(c[20]), .CI(n239), .CON(n286), 
        .SN(n285) );
  AND2x2_ASAP7_6t_L U84 ( .A(p[8]), .B(p[1]), .Y(n19) );
  AND2x2_ASAP7_6t_L U85 ( .A(s[11]), .B(n258), .Y(n20) );
  XOR2xp5r_ASAP7_6t_L U86 ( .A(p[1]), .B(p[8]), .Y(out[1]) );
  XOR2xp5r_ASAP7_6t_L U87 ( .A(n258), .B(s[11]), .Y(out[4]) );
  XOR2xp5r_ASAP7_6t_L U88 ( .A(n253), .B(n237), .Y(out[15]) );
  XOR2xp5r_ASAP7_6t_L U89 ( .A(n24), .B(n25), .Y(s[9]) );
  NAND2xp5R_ASAP7_6t_L U90 ( .A(b[1]), .B(a[1]), .Y(n24) );
  XOR2xp5r_ASAP7_6t_L U91 ( .A(n26), .B(n27), .Y(s[21]) );
  XOR2xp5r_ASAP7_6t_L U92 ( .A(n28), .B(n29), .Y(s[20]) );
  XOR2xp5r_ASAP7_6t_L U93 ( .A(n30), .B(n31), .Y(s[19]) );
  XOR2xp5r_ASAP7_6t_L U94 ( .A(n32), .B(n33), .Y(s[18]) );
  XOR2xp5r_ASAP7_6t_L U95 ( .A(n34), .B(n35), .Y(s[17]) );
  XOR2xp5r_ASAP7_6t_L U96 ( .A(n36), .B(n37), .Y(s[16]) );
  XOR2xp5r_ASAP7_6t_L U97 ( .A(n38), .B(n39), .Y(s[15]) );
  XOR2xp5r_ASAP7_6t_L U98 ( .A(n40), .B(n41), .Y(s[14]) );
  XOR2xp5r_ASAP7_6t_L U99 ( .A(n42), .B(n43), .Y(s[13]) );
  XOR2xp5r_ASAP7_6t_L U100 ( .A(n44), .B(n45), .Y(s[12]) );
  XOR2xp5r_ASAP7_6t_L U101 ( .A(n46), .B(n47), .Y(s[11]) );
  NOR2xp5_ASAP7_6t_L U102 ( .A(n48), .B(n49), .Y(p[8]) );
  NOR2xp5_ASAP7_6t_L U103 ( .A(n50), .B(n51), .Y(p[1]) );
  NOR2xp5_ASAP7_6t_L U104 ( .A(n52), .B(n49), .Y(p[16]) );
  NOR2xp5_ASAP7_6t_L U105 ( .A(n50), .B(n49), .Y(out[0]) );
  INVx1_ASAP7_6t_L U106 ( .A(n286), .Y(n237) );
  INVx1_ASAP7_6t_L U107 ( .A(n285), .Y(out[14]) );
  INVx1_ASAP7_6t_L U108 ( .A(n284), .Y(n239) );
  INVx1_ASAP7_6t_L U109 ( .A(n283), .Y(out[13]) );
  INVx1_ASAP7_6t_L U110 ( .A(n282), .Y(n241) );
  INVx1_ASAP7_6t_L U111 ( .A(n281), .Y(out[12]) );
  INVx1_ASAP7_6t_L U112 ( .A(n280), .Y(n243) );
  INVx1_ASAP7_6t_L U113 ( .A(n279), .Y(out[11]) );
  INVx1_ASAP7_6t_L U114 ( .A(n278), .Y(n245) );
  INVx1_ASAP7_6t_L U115 ( .A(n277), .Y(out[10]) );
  INVx1_ASAP7_6t_L U116 ( .A(n276), .Y(n247) );
  INVx1_ASAP7_6t_L U117 ( .A(n275), .Y(out[9]) );
  INVx1_ASAP7_6t_L U118 ( .A(n274), .Y(n249) );
  INVx1_ASAP7_6t_L U119 ( .A(n273), .Y(out[8]) );
  INVx1_ASAP7_6t_L U120 ( .A(n272), .Y(n251) );
  INVx1_ASAP7_6t_L U121 ( .A(n271), .Y(out[7]) );
  OAI22xp5_ASAP7_6t_L U122 ( .A1(n27), .A2(n26), .B1(n53), .B2(n54), .Y(n253)
         );
  OAI211xp33_ASAP7_6t_L U123 ( .A1(n53), .A2(n54), .B(b[7]), .C(a[7]), .Y(n27)
         );
  INVx1_ASAP7_6t_L U124 ( .A(n270), .Y(n254) );
  INVx1_ASAP7_6t_L U125 ( .A(n269), .Y(out[6]) );
  INVx1_ASAP7_6t_L U126 ( .A(n268), .Y(n256) );
  INVx1_ASAP7_6t_L U127 ( .A(n267), .Y(out[5]) );
  INVx1_ASAP7_6t_L U128 ( .A(n266), .Y(n258) );
  INVx1_ASAP7_6t_L U129 ( .A(n265), .Y(out[3]) );
  INVx1_ASAP7_6t_L U130 ( .A(n264), .Y(n261) );
  INVx1_ASAP7_6t_L U131 ( .A(n263), .Y(out[2]) );
  NOR3x1f_ASAP7_6t_L U132 ( .A(n25), .B(n48), .C(n51), .Y(c[9]) );
  NAND2xp5R_ASAP7_6t_L U133 ( .A(b[2]), .B(a[0]), .Y(n25) );
  NOR2xp5_ASAP7_6t_L U134 ( .A(n29), .B(n28), .Y(c[20]) );
  OAI21xp25_ASAP7_6t_L U135 ( .A1(n54), .A2(n55), .B(n26), .Y(n28) );
  NAND2xp5R_ASAP7_6t_L U136 ( .A(n54), .B(n55), .Y(n26) );
  OAI21xp25_ASAP7_6t_L U137 ( .A1(n56), .A2(n57), .B(n58), .Y(n55) );
  XOR2xp5r_ASAP7_6t_L U138 ( .A(n59), .B(n53), .Y(n54) );
  NAND2xp5R_ASAP7_6t_L U139 ( .A(a[6]), .B(b[7]), .Y(n53) );
  NAND2xp5R_ASAP7_6t_L U140 ( .A(b[6]), .B(a[7]), .Y(n59) );
  NOR2xp5_ASAP7_6t_L U141 ( .A(n31), .B(n30), .Y(c[19]) );
  OAI21xp25_ASAP7_6t_L U142 ( .A1(n60), .A2(n61), .B(n29), .Y(n30) );
  NAND2xp5R_ASAP7_6t_L U143 ( .A(n60), .B(n61), .Y(n29) );
  OR2x2_ASAP7_6t_L U144 ( .A(n62), .B(n63), .Y(n61) );
  NOR3x1f_ASAP7_6t_L U145 ( .A(n64), .B(n65), .C(n66), .Y(n63) );
  NOR3x1f_ASAP7_6t_L U146 ( .A(n67), .B(n68), .C(n69), .Y(n62) );
  INVx1_ASAP7_6t_L U147 ( .A(n64), .Y(n67) );
  INVx1_ASAP7_6t_L U148 ( .A(n70), .Y(n60) );
  A2O1A1Ixp33_ASAP7_6t_L U149 ( .A1(b[5]), .A2(a[7]), .B(n57), .C(n58), .Y(n70) );
  NAND3xp33R_ASAP7_6t_L U150 ( .A(b[5]), .B(n57), .C(a[7]), .Y(n58) );
  XOR2xp5r_ASAP7_6t_L U151 ( .A(n71), .B(n56), .Y(n57) );
  NAND2xp5R_ASAP7_6t_L U152 ( .A(b[7]), .B(a[5]), .Y(n56) );
  NAND2xp5R_ASAP7_6t_L U153 ( .A(a[6]), .B(b[6]), .Y(n71) );
  OA22x1_ASAP7_6t_L U154 ( .A1(n72), .A2(n73), .B1(n74), .B2(n75), .Y(n31) );
  AO21x1_ASAP7_6t_L U155 ( .A1(n32), .A2(n33), .B(n76), .Y(c[18]) );
  NOR3x1f_ASAP7_6t_L U156 ( .A(n33), .B(n77), .C(n78), .Y(n76) );
  XOR2xp5r_ASAP7_6t_L U157 ( .A(n79), .B(n75), .Y(n33) );
  AOI21xp25_ASAP7_6t_L U158 ( .A1(n80), .A2(n81), .B(n82), .Y(n75) );
  NOR3x1f_ASAP7_6t_L U159 ( .A(n81), .B(n83), .C(n78), .Y(n82) );
  XOR2xp5r_ASAP7_6t_L U160 ( .A(n84), .B(n74), .Y(n79) );
  INVx1_ASAP7_6t_L U161 ( .A(n72), .Y(n74) );
  XOR2xp5r_ASAP7_6t_L U162 ( .A(n85), .B(n64), .Y(n72) );
  XOR2xp5r_ASAP7_6t_L U163 ( .A(n86), .B(n87), .Y(n64) );
  NAND2xp5R_ASAP7_6t_L U164 ( .A(a[4]), .B(b[7]), .Y(n87) );
  AOI22xp25_ASAP7_6t_L U165 ( .A1(n88), .A2(n89), .B1(n90), .B2(n91), .Y(n86)
         );
  XOR2xp5r_ASAP7_6t_L U166 ( .A(n92), .B(n73), .Y(n85) );
  NAND2xp5R_ASAP7_6t_L U167 ( .A(b[5]), .B(a[6]), .Y(n73) );
  NAND2xp5R_ASAP7_6t_L U168 ( .A(b[6]), .B(a[5]), .Y(n92) );
  NOR2xp5_ASAP7_6t_L U169 ( .A(n77), .B(n78), .Y(n84) );
  OAI22xp5_ASAP7_6t_L U170 ( .A1(n93), .A2(n94), .B1(n95), .B2(n96), .Y(n32)
         );
  INVx1_ASAP7_6t_L U171 ( .A(n97), .Y(n95) );
  AO21x1_ASAP7_6t_L U172 ( .A1(n34), .A2(n35), .B(n98), .Y(c[17]) );
  NOR3x1f_ASAP7_6t_L U173 ( .A(n34), .B(n77), .C(n99), .Y(n98) );
  OAI22xp5_ASAP7_6t_L U174 ( .A1(n100), .A2(n101), .B1(n102), .B2(n103), .Y(
        n35) );
  INVx1_ASAP7_6t_L U175 ( .A(n101), .Y(n102) );
  XOR2xp5r_ASAP7_6t_L U176 ( .A(n104), .B(n93), .Y(n34) );
  AOI22xp25_ASAP7_6t_L U177 ( .A1(n105), .A2(n106), .B1(n107), .B2(n108), .Y(
        n93) );
  XOR2xp5r_ASAP7_6t_L U178 ( .A(n109), .B(n94), .Y(n104) );
  INVx1_ASAP7_6t_L U179 ( .A(n96), .Y(n94) );
  XOR2xp5r_ASAP7_6t_L U180 ( .A(n81), .B(n110), .Y(n96) );
  XOR2xp5r_ASAP7_6t_L U181 ( .A(n97), .B(n111), .Y(n110) );
  NAND2xp5R_ASAP7_6t_L U182 ( .A(b[4]), .B(a[6]), .Y(n111) );
  OAI22xp5_ASAP7_6t_L U183 ( .A1(n112), .A2(n113), .B1(n114), .B2(n115), .Y(
        n97) );
  XOR2xp5r_ASAP7_6t_L U184 ( .A(n116), .B(n80), .Y(n81) );
  XOR2xp5r_ASAP7_6t_L U185 ( .A(n91), .B(n90), .Y(n80) );
  AND2x2_ASAP7_6t_L U186 ( .A(b[5]), .B(a[5]), .Y(n90) );
  XOR2xp5r_ASAP7_6t_L U187 ( .A(n89), .B(n88), .Y(n91) );
  NOR2xp5_ASAP7_6t_L U188 ( .A(n66), .B(n69), .Y(n88) );
  NOR2xp5_ASAP7_6t_L U189 ( .A(n117), .B(n65), .Y(n89) );
  AOI22xp25_ASAP7_6t_L U190 ( .A1(n118), .A2(n119), .B1(n120), .B2(n121), .Y(
        n116) );
  NOR2xp5_ASAP7_6t_L U191 ( .A(n77), .B(n99), .Y(n109) );
  OAI22xp5_ASAP7_6t_L U192 ( .A1(n36), .A2(n37), .B1(n122), .B2(n123), .Y(
        c[16]) );
  INVx1_ASAP7_6t_L U193 ( .A(n37), .Y(n122) );
  XOR2xp5r_ASAP7_6t_L U194 ( .A(n123), .B(n124), .Y(n37) );
  XOR2xp5r_ASAP7_6t_L U195 ( .A(n100), .B(n101), .Y(n124) );
  XOR2xp5r_ASAP7_6t_L U196 ( .A(n103), .B(n125), .Y(n101) );
  XOR2xp5r_ASAP7_6t_L U197 ( .A(n106), .B(n105), .Y(n125) );
  INVx1_ASAP7_6t_L U198 ( .A(n107), .Y(n105) );
  XOR2xp5r_ASAP7_6t_L U199 ( .A(n126), .B(n108), .Y(n107) );
  XOR2xp5r_ASAP7_6t_L U200 ( .A(n121), .B(n120), .Y(n108) );
  AND2x2_ASAP7_6t_L U201 ( .A(a[4]), .B(b[5]), .Y(n120) );
  XOR2xp5r_ASAP7_6t_L U202 ( .A(n118), .B(n119), .Y(n121) );
  NOR2xp5_ASAP7_6t_L U203 ( .A(n52), .B(n65), .Y(n119) );
  INVx1_ASAP7_6t_L U204 ( .A(b[7]), .Y(n65) );
  NOR2xp5_ASAP7_6t_L U205 ( .A(n117), .B(n69), .Y(n118) );
  AOI21xp25_ASAP7_6t_L U206 ( .A1(n127), .A2(n128), .B(n129), .Y(n126) );
  NOR3x1f_ASAP7_6t_L U207 ( .A(n128), .B(n68), .C(n99), .Y(n129) );
  XOR2xp5r_ASAP7_6t_L U208 ( .A(n112), .B(n113), .Y(n106) );
  NAND2xp5R_ASAP7_6t_L U209 ( .A(a[7]), .B(b[2]), .Y(n113) );
  XOR2xp5r_ASAP7_6t_L U210 ( .A(n130), .B(n114), .Y(n112) );
  NAND2xp5R_ASAP7_6t_L U211 ( .A(b[4]), .B(a[5]), .Y(n114) );
  INVx1_ASAP7_6t_L U212 ( .A(n115), .Y(n130) );
  NAND2xp5R_ASAP7_6t_L U213 ( .A(b[3]), .B(a[6]), .Y(n115) );
  OA22x1_ASAP7_6t_L U214 ( .A1(n131), .A2(n132), .B1(n133), .B2(n134), .Y(n103) );
  INVx1_ASAP7_6t_L U215 ( .A(n131), .Y(n133) );
  AOI21xp25_ASAP7_6t_L U216 ( .A1(n135), .A2(n136), .B(n137), .Y(n100) );
  NOR3x1f_ASAP7_6t_L U217 ( .A(n136), .B(n138), .C(n83), .Y(n137) );
  AOI21xp25_ASAP7_6t_L U218 ( .A1(n139), .A2(n140), .B(n141), .Y(n123) );
  NOR3x1f_ASAP7_6t_L U219 ( .A(n139), .B(n66), .C(n78), .Y(n141) );
  AOI22xp25_ASAP7_6t_L U220 ( .A1(n142), .A2(n143), .B1(n144), .B2(n145), .Y(
        n36) );
  AO21x1_ASAP7_6t_L U221 ( .A1(n39), .A2(n38), .B(n146), .Y(c[15]) );
  NOR3x1f_ASAP7_6t_L U222 ( .A(n39), .B(n51), .C(n77), .Y(n146) );
  OAI22xp5_ASAP7_6t_L U223 ( .A1(n147), .A2(n148), .B1(n149), .B2(n150), .Y(
        n38) );
  INVx1_ASAP7_6t_L U224 ( .A(n151), .Y(n148) );
  XOR2xp5r_ASAP7_6t_L U225 ( .A(n142), .B(n152), .Y(n39) );
  XOR2xp5r_ASAP7_6t_L U226 ( .A(n153), .B(n143), .Y(n152) );
  INVx1_ASAP7_6t_L U227 ( .A(n144), .Y(n143) );
  XOR2xp5r_ASAP7_6t_L U228 ( .A(n154), .B(n136), .Y(n144) );
  XOR2xp5r_ASAP7_6t_L U229 ( .A(n155), .B(n135), .Y(n136) );
  XOR2xp5r_ASAP7_6t_L U230 ( .A(n127), .B(n128), .Y(n135) );
  XOR2xp5r_ASAP7_6t_L U231 ( .A(n156), .B(n140), .Y(n128) );
  OAI22xp5_ASAP7_6t_L U232 ( .A1(n157), .A2(n158), .B1(n159), .B2(n160), .Y(
        n140) );
  INVx1_ASAP7_6t_L U233 ( .A(n157), .Y(n159) );
  XOR2xp5r_ASAP7_6t_L U234 ( .A(n161), .B(n139), .Y(n156) );
  XOR2xp5r_ASAP7_6t_L U235 ( .A(n131), .B(n162), .Y(n139) );
  XOR2xp5r_ASAP7_6t_L U236 ( .A(n163), .B(n132), .Y(n162) );
  NAND2xp5R_ASAP7_6t_L U237 ( .A(a[3]), .B(b[5]), .Y(n132) );
  NOR2xp5_ASAP7_6t_L U238 ( .A(n66), .B(n78), .Y(n163) );
  XOR2xp5r_ASAP7_6t_L U239 ( .A(n164), .B(n134), .Y(n131) );
  NAND2xp5R_ASAP7_6t_L U240 ( .A(b[7]), .B(a[1]), .Y(n134) );
  NOR2xp5_ASAP7_6t_L U241 ( .A(n69), .B(n52), .Y(n164) );
  NOR2xp5_ASAP7_6t_L U242 ( .A(n68), .B(n99), .Y(n161) );
  NOR3x1f_ASAP7_6t_L U243 ( .A(n165), .B(n117), .C(n78), .Y(n127) );
  INVx1_ASAP7_6t_L U244 ( .A(n166), .Y(n165) );
  NAND2xp5R_ASAP7_6t_L U245 ( .A(n167), .B(n168), .Y(n155) );
  NOR3x1f_ASAP7_6t_L U246 ( .A(n83), .B(n145), .C(n138), .Y(n154) );
  NOR3x1f_ASAP7_6t_L U247 ( .A(n169), .B(n51), .C(n83), .Y(n145) );
  NOR2xp5_ASAP7_6t_L U248 ( .A(n51), .B(n77), .Y(n153) );
  OAI22xp5_ASAP7_6t_L U249 ( .A1(n170), .A2(n168), .B1(n171), .B2(n172), .Y(
        n142) );
  INVx1_ASAP7_6t_L U250 ( .A(n170), .Y(n171) );
  AO21x1_ASAP7_6t_L U251 ( .A1(n40), .A2(n41), .B(n173), .Y(c[14]) );
  NOR3x1f_ASAP7_6t_L U252 ( .A(n41), .B(n77), .C(n49), .Y(n173) );
  XOR2xp5r_ASAP7_6t_L U253 ( .A(n174), .B(n175), .Y(n41) );
  XOR2xp5r_ASAP7_6t_L U254 ( .A(n176), .B(n147), .Y(n175) );
  INVx1_ASAP7_6t_L U255 ( .A(n149), .Y(n147) );
  XOR2xp5r_ASAP7_6t_L U256 ( .A(n172), .B(n177), .Y(n149) );
  XOR2xp5r_ASAP7_6t_L U257 ( .A(n151), .B(n170), .Y(n177) );
  XOR2xp5r_ASAP7_6t_L U258 ( .A(n178), .B(n168), .Y(n170) );
  XOR2xp5r_ASAP7_6t_L U259 ( .A(n166), .B(n167), .Y(n168) );
  NOR2xp5_ASAP7_6t_L U260 ( .A(n99), .B(n66), .Y(n167) );
  XOR2xp5r_ASAP7_6t_L U261 ( .A(n179), .B(n157), .Y(n166) );
  XOR2xp5r_ASAP7_6t_L U262 ( .A(n180), .B(n160), .Y(n157) );
  NAND2xp5R_ASAP7_6t_L U263 ( .A(b[7]), .B(a[0]), .Y(n160) );
  NOR2xp5_ASAP7_6t_L U264 ( .A(n48), .B(n69), .Y(n180) );
  INVx1_ASAP7_6t_L U265 ( .A(a[1]), .Y(n48) );
  XOR2xp5r_ASAP7_6t_L U266 ( .A(n181), .B(n158), .Y(n179) );
  NAND2xp5R_ASAP7_6t_L U267 ( .A(a[2]), .B(b[5]), .Y(n158) );
  NAND2xp5R_ASAP7_6t_L U268 ( .A(b[4]), .B(a[3]), .Y(n181) );
  AOI22xp25_ASAP7_6t_L U269 ( .A1(n182), .A2(n183), .B1(n184), .B2(n185), .Y(
        n178) );
  NOR3x1f_ASAP7_6t_L U270 ( .A(n186), .B(n138), .C(n66), .Y(n151) );
  XOR2xp5r_ASAP7_6t_L U271 ( .A(n187), .B(n169), .Y(n172) );
  NAND2xp5R_ASAP7_6t_L U272 ( .A(a[5]), .B(b[2]), .Y(n169) );
  NOR2xp5_ASAP7_6t_L U273 ( .A(n51), .B(n83), .Y(n187) );
  NOR2xp5_ASAP7_6t_L U274 ( .A(n77), .B(n49), .Y(n176) );
  INVx1_ASAP7_6t_L U275 ( .A(a[7]), .Y(n77) );
  INVx1_ASAP7_6t_L U276 ( .A(n150), .Y(n174) );
  AOI22xp25_ASAP7_6t_L U277 ( .A1(n188), .A2(n189), .B1(n190), .B2(n191), .Y(
        n150) );
  INVx1_ASAP7_6t_L U278 ( .A(n188), .Y(n190) );
  AO21x1_ASAP7_6t_L U279 ( .A1(n192), .A2(n193), .B(n194), .Y(n40) );
  NOR3x1f_ASAP7_6t_L U280 ( .A(n192), .B(n51), .C(n68), .Y(n194) );
  AO21x1_ASAP7_6t_L U281 ( .A1(n43), .A2(n42), .B(n195), .Y(c[13]) );
  NOR3x1f_ASAP7_6t_L U282 ( .A(n43), .B(n83), .C(n49), .Y(n195) );
  OAI22xp5_ASAP7_6t_L U283 ( .A1(n196), .A2(n197), .B1(n198), .B2(n199), .Y(
        n42) );
  INVx1_ASAP7_6t_L U284 ( .A(n197), .Y(n198) );
  XOR2xp5r_ASAP7_6t_L U285 ( .A(n193), .B(n200), .Y(n43) );
  XOR2xp5r_ASAP7_6t_L U286 ( .A(n201), .B(n192), .Y(n200) );
  XOR2xp5r_ASAP7_6t_L U287 ( .A(n202), .B(n188), .Y(n192) );
  XOR2xp5r_ASAP7_6t_L U288 ( .A(n203), .B(n191), .Y(n188) );
  XOR2xp5r_ASAP7_6t_L U289 ( .A(n185), .B(n184), .Y(n191) );
  NOR2xp5_ASAP7_6t_L U290 ( .A(n78), .B(n52), .Y(n184) );
  XOR2xp5r_ASAP7_6t_L U291 ( .A(n182), .B(n183), .Y(n185) );
  NOR2xp5_ASAP7_6t_L U292 ( .A(n69), .B(n50), .Y(n183) );
  INVx1_ASAP7_6t_L U293 ( .A(b[6]), .Y(n69) );
  AND2x2_ASAP7_6t_L U294 ( .A(b[5]), .B(a[1]), .Y(n182) );
  NOR2xp5_ASAP7_6t_L U295 ( .A(n204), .B(n205), .Y(n203) );
  XOR2xp5r_ASAP7_6t_L U296 ( .A(n206), .B(n189), .Y(n202) );
  XOR2xp5r_ASAP7_6t_L U297 ( .A(n207), .B(n186), .Y(n189) );
  NAND2xp5R_ASAP7_6t_L U298 ( .A(b[3]), .B(a[3]), .Y(n186) );
  NAND2xp5R_ASAP7_6t_L U299 ( .A(b[2]), .B(a[4]), .Y(n207) );
  NOR2xp5_ASAP7_6t_L U300 ( .A(n51), .B(n68), .Y(n206) );
  NOR2xp5_ASAP7_6t_L U301 ( .A(n83), .B(n49), .Y(n201) );
  INVx1_ASAP7_6t_L U302 ( .A(a[6]), .Y(n83) );
  AO21x1_ASAP7_6t_L U303 ( .A1(n208), .A2(n209), .B(n210), .Y(n193) );
  NOR3x1f_ASAP7_6t_L U304 ( .A(n209), .B(n138), .C(n117), .Y(n210) );
  INVx1_ASAP7_6t_L U305 ( .A(a[3]), .Y(n117) );
  AO21x1_ASAP7_6t_L U306 ( .A1(n44), .A2(n45), .B(n211), .Y(c[12]) );
  NOR3x1f_ASAP7_6t_L U307 ( .A(n44), .B(n68), .C(n49), .Y(n211) );
  OAI22xp5_ASAP7_6t_L U308 ( .A1(n212), .A2(n213), .B1(n214), .B2(n215), .Y(
        n45) );
  XOR2xp5r_ASAP7_6t_L U309 ( .A(n196), .B(n216), .Y(n44) );
  XOR2xp5r_ASAP7_6t_L U310 ( .A(n217), .B(n197), .Y(n216) );
  XOR2xp5r_ASAP7_6t_L U311 ( .A(n218), .B(n209), .Y(n197) );
  XOR2xp5r_ASAP7_6t_L U312 ( .A(n208), .B(n219), .Y(n209) );
  NAND2xp5R_ASAP7_6t_L U313 ( .A(b[3]), .B(a[2]), .Y(n219) );
  XOR2xp5r_ASAP7_6t_L U314 ( .A(n205), .B(n204), .Y(n208) );
  NAND2xp5R_ASAP7_6t_L U315 ( .A(b[4]), .B(a[1]), .Y(n204) );
  NAND2xp5R_ASAP7_6t_L U316 ( .A(b[5]), .B(a[0]), .Y(n205) );
  XOR2xp5r_ASAP7_6t_L U317 ( .A(n220), .B(n199), .Y(n218) );
  NAND2xp5R_ASAP7_6t_L U318 ( .A(a[4]), .B(b[1]), .Y(n199) );
  NAND2xp5R_ASAP7_6t_L U319 ( .A(a[3]), .B(b[2]), .Y(n220) );
  NOR2xp5_ASAP7_6t_L U320 ( .A(n68), .B(n49), .Y(n217) );
  INVx1_ASAP7_6t_L U321 ( .A(a[5]), .Y(n68) );
  AOI21xp25_ASAP7_6t_L U322 ( .A1(n221), .A2(n222), .B(n223), .Y(n196) );
  NOR3x1f_ASAP7_6t_L U323 ( .A(n222), .B(n138), .C(n52), .Y(n223) );
  AO21x1_ASAP7_6t_L U324 ( .A1(n46), .A2(n47), .B(n224), .Y(c[11]) );
  NOR3x1f_ASAP7_6t_L U325 ( .A(n47), .B(n66), .C(n49), .Y(n224) );
  XOR2xp5r_ASAP7_6t_L U326 ( .A(n225), .B(n212), .Y(n47) );
  AOI21xp25_ASAP7_6t_L U327 ( .A1(n226), .A2(n227), .B(n228), .Y(n212) );
  NOR3x1f_ASAP7_6t_L U328 ( .A(n227), .B(n51), .C(n52), .Y(n228) );
  XOR2xp5r_ASAP7_6t_L U329 ( .A(n229), .B(n213), .Y(n225) );
  INVx1_ASAP7_6t_L U330 ( .A(n214), .Y(n213) );
  XOR2xp5r_ASAP7_6t_L U331 ( .A(n222), .B(n230), .Y(n214) );
  XOR2xp5r_ASAP7_6t_L U332 ( .A(n231), .B(n215), .Y(n230) );
  NAND2xp5R_ASAP7_6t_L U333 ( .A(a[3]), .B(b[1]), .Y(n215) );
  NOR2xp5_ASAP7_6t_L U334 ( .A(n138), .B(n52), .Y(n231) );
  INVx1_ASAP7_6t_L U335 ( .A(b[2]), .Y(n138) );
  XOR2xp5r_ASAP7_6t_L U336 ( .A(n232), .B(n221), .Y(n222) );
  NOR2xp5_ASAP7_6t_L U337 ( .A(n78), .B(n50), .Y(n221) );
  INVx1_ASAP7_6t_L U338 ( .A(b[4]), .Y(n78) );
  NAND2xp5R_ASAP7_6t_L U339 ( .A(a[1]), .B(b[3]), .Y(n232) );
  NOR2xp5_ASAP7_6t_L U340 ( .A(n66), .B(n49), .Y(n229) );
  INVx1_ASAP7_6t_L U341 ( .A(b[0]), .Y(n49) );
  INVx1_ASAP7_6t_L U342 ( .A(a[4]), .Y(n66) );
  NOR2xp5_ASAP7_6t_L U343 ( .A(n233), .B(n260), .Y(n46) );
  XOR2xp5r_ASAP7_6t_L U344 ( .A(n227), .B(n234), .Y(n260) );
  XOR2xp5r_ASAP7_6t_L U345 ( .A(n235), .B(n233), .Y(n234) );
  NOR2xp5_ASAP7_6t_L U346 ( .A(n51), .B(n52), .Y(n235) );
  INVx1_ASAP7_6t_L U347 ( .A(a[2]), .Y(n52) );
  INVx1_ASAP7_6t_L U348 ( .A(b[1]), .Y(n51) );
  XOR2xp5r_ASAP7_6t_L U349 ( .A(n236), .B(n226), .Y(n227) );
  NOR2xp5_ASAP7_6t_L U350 ( .A(n99), .B(n50), .Y(n226) );
  INVx1_ASAP7_6t_L U351 ( .A(a[0]), .Y(n50) );
  INVx1_ASAP7_6t_L U352 ( .A(b[3]), .Y(n99) );
  NAND2xp5R_ASAP7_6t_L U353 ( .A(b[2]), .B(a[1]), .Y(n236) );
  NAND2xp5R_ASAP7_6t_L U354 ( .A(b[0]), .B(a[3]), .Y(n233) );
endmodule

