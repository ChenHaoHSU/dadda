
module DADDA_8x8 ( a, b, out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] out;
  wire   c_30_, add_98_CI, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n225, n227, n229, n231, n233, n235, n237, n239, n240,
         n241, n242, n243, n244, n245, n246, n248, n249, n251, n252, n254,
         n255, n257, n258, n260, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289;
  wire   [63:1] p;
  wire   [41:30] s;

  FAxp33_ASAP7_6t_L add_98_U1_0 ( .A(p[1]), .B(p[8]), .CI(add_98_CI), .CON(
        n263), .SN(n262) );
  FAxp33_ASAP7_6t_L add_98_U1_1 ( .A(s[30]), .B(p[16]), .CI(n260), .CON(n265), 
        .SN(n264) );
  FAxp33_ASAP7_6t_L add_98_U1_2 ( .A(c_30_), .B(s[31]), .CI(n258), .CON(n267), 
        .SN(n266) );
  FAxp33_ASAP7_6t_L add_98_U1_3 ( .A(n257), .B(s[32]), .CI(n255), .CON(n269), 
        .SN(n268) );
  FAxp33_ASAP7_6t_L add_98_U1_4 ( .A(n254), .B(s[33]), .CI(n252), .CON(n271), 
        .SN(n270) );
  FAxp33_ASAP7_6t_L add_98_U1_5 ( .A(n251), .B(s[34]), .CI(n249), .CON(n273), 
        .SN(n272) );
  FAxp33_ASAP7_6t_L add_98_U1_6 ( .A(n248), .B(s[35]), .CI(n246), .CON(n275), 
        .SN(n274) );
  FAxp33_ASAP7_6t_L add_98_U1_7 ( .A(n239), .B(s[36]), .CI(n237), .CON(n277), 
        .SN(n276) );
  FAxp33_ASAP7_6t_L add_98_U1_8 ( .A(n241), .B(s[37]), .CI(n235), .CON(n279), 
        .SN(n278) );
  FAxp33_ASAP7_6t_L add_98_U1_9 ( .A(n240), .B(s[38]), .CI(n233), .CON(n281), 
        .SN(n280) );
  FAxp33_ASAP7_6t_L add_98_U1_10 ( .A(n242), .B(s[39]), .CI(n231), .CON(n283), 
        .SN(n282) );
  FAxp33_ASAP7_6t_L add_98_U1_11 ( .A(n243), .B(s[40]), .CI(n229), .CON(n285), 
        .SN(n284) );
  FAxp33_ASAP7_6t_L add_98_U1_12 ( .A(n244), .B(s[41]), .CI(n227), .CON(n287), 
        .SN(n286) );
  FAxp33_ASAP7_6t_L add_98_U1_13 ( .A(n245), .B(p[63]), .CI(n225), .CON(n289), 
        .SN(n288) );
  TIELOxp5_ASAP7_6t_L U83 ( .L(add_98_CI) );
  XOR2xp5r_ASAP7_6t_L U84 ( .A(n19), .B(n20), .Y(s[41]) );
  NAND2xp5R_ASAP7_6t_L U85 ( .A(a[7]), .B(b[6]), .Y(n19) );
  XOR2xp5r_ASAP7_6t_L U86 ( .A(n21), .B(n22), .Y(s[40]) );
  NOR2xp5_ASAP7_6t_L U87 ( .A(n23), .B(n24), .Y(n21) );
  XOR2xp5r_ASAP7_6t_L U88 ( .A(n25), .B(n26), .Y(s[39]) );
  NOR2xp5_ASAP7_6t_L U89 ( .A(n23), .B(n27), .Y(n25) );
  XOR2xp5r_ASAP7_6t_L U90 ( .A(n28), .B(n29), .Y(s[38]) );
  XOR2xp5r_ASAP7_6t_L U91 ( .A(n30), .B(n31), .Y(s[37]) );
  XOR2xp5r_ASAP7_6t_L U92 ( .A(n32), .B(n33), .Y(s[36]) );
  XOR2xp5r_ASAP7_6t_L U93 ( .A(n34), .B(n35), .Y(s[35]) );
  XOR2xp5r_ASAP7_6t_L U94 ( .A(n36), .B(n37), .Y(s[34]) );
  XOR2xp5r_ASAP7_6t_L U95 ( .A(n38), .B(n39), .Y(s[33]) );
  NAND2xp5R_ASAP7_6t_L U96 ( .A(a[5]), .B(b[0]), .Y(n38) );
  XOR2xp5r_ASAP7_6t_L U97 ( .A(n40), .B(n41), .Y(s[32]) );
  NOR2xp5_ASAP7_6t_L U98 ( .A(n42), .B(n43), .Y(n40) );
  XOR2xp5r_ASAP7_6t_L U99 ( .A(n44), .B(n45), .Y(s[31]) );
  NOR2xp5_ASAP7_6t_L U100 ( .A(n46), .B(n43), .Y(n44) );
  XOR2xp5r_ASAP7_6t_L U101 ( .A(n47), .B(n48), .Y(s[30]) );
  NAND2xp5R_ASAP7_6t_L U102 ( .A(b[1]), .B(a[1]), .Y(n47) );
  NOR2xp5_ASAP7_6t_L U103 ( .A(n49), .B(n43), .Y(p[8]) );
  NOR2xp5_ASAP7_6t_L U104 ( .A(n23), .B(n50), .Y(p[63]) );
  NOR2xp5_ASAP7_6t_L U105 ( .A(n51), .B(n52), .Y(p[1]) );
  NOR2xp5_ASAP7_6t_L U106 ( .A(n53), .B(n43), .Y(p[16]) );
  NOR2xp5_ASAP7_6t_L U107 ( .A(n52), .B(n43), .Y(out[0]) );
  INVx1_ASAP7_6t_L U108 ( .A(n289), .Y(out[15]) );
  INVx1_ASAP7_6t_L U109 ( .A(n288), .Y(out[14]) );
  INVx1_ASAP7_6t_L U110 ( .A(n287), .Y(n225) );
  INVx1_ASAP7_6t_L U111 ( .A(n286), .Y(out[13]) );
  INVx1_ASAP7_6t_L U112 ( .A(n285), .Y(n227) );
  INVx1_ASAP7_6t_L U113 ( .A(n284), .Y(out[12]) );
  INVx1_ASAP7_6t_L U114 ( .A(n283), .Y(n229) );
  INVx1_ASAP7_6t_L U115 ( .A(n282), .Y(out[11]) );
  INVx1_ASAP7_6t_L U116 ( .A(n281), .Y(n231) );
  INVx1_ASAP7_6t_L U117 ( .A(n280), .Y(out[10]) );
  INVx1_ASAP7_6t_L U118 ( .A(n279), .Y(n233) );
  INVx1_ASAP7_6t_L U119 ( .A(n278), .Y(out[9]) );
  INVx1_ASAP7_6t_L U120 ( .A(n277), .Y(n235) );
  INVx1_ASAP7_6t_L U121 ( .A(n276), .Y(out[8]) );
  INVx1_ASAP7_6t_L U122 ( .A(n275), .Y(n237) );
  INVx1_ASAP7_6t_L U123 ( .A(n274), .Y(out[7]) );
  OAI22xp5_ASAP7_6t_L U124 ( .A1(n54), .A2(n55), .B1(n34), .B2(n35), .Y(n239)
         );
  XOR2xp5r_ASAP7_6t_L U125 ( .A(n56), .B(n55), .Y(n35) );
  INVx1_ASAP7_6t_L U126 ( .A(n54), .Y(n56) );
  XOR2xp5r_ASAP7_6t_L U127 ( .A(n57), .B(n58), .Y(n34) );
  INVx1_ASAP7_6t_L U128 ( .A(n59), .Y(n57) );
  XOR2xp5r_ASAP7_6t_L U129 ( .A(n60), .B(n61), .Y(n55) );
  AOI22xp25_ASAP7_6t_L U130 ( .A1(n62), .A2(n63), .B1(n64), .B2(n65), .Y(n54)
         );
  OAI22xp5_ASAP7_6t_L U131 ( .A1(n66), .A2(n67), .B1(n30), .B2(n31), .Y(n240)
         );
  XOR2xp5r_ASAP7_6t_L U132 ( .A(n68), .B(n67), .Y(n31) );
  INVx1_ASAP7_6t_L U133 ( .A(n66), .Y(n68) );
  XOR2xp5r_ASAP7_6t_L U134 ( .A(n69), .B(n70), .Y(n30) );
  INVx1_ASAP7_6t_L U135 ( .A(n71), .Y(n69) );
  XOR2xp5r_ASAP7_6t_L U136 ( .A(n72), .B(n73), .Y(n67) );
  AOI22xp25_ASAP7_6t_L U137 ( .A1(n74), .A2(n75), .B1(n76), .B2(n77), .Y(n66)
         );
  OAI22xp5_ASAP7_6t_L U138 ( .A1(n78), .A2(n79), .B1(n32), .B2(n33), .Y(n241)
         );
  XOR2xp5r_ASAP7_6t_L U139 ( .A(n78), .B(n80), .Y(n33) );
  XOR2xp5r_ASAP7_6t_L U140 ( .A(n81), .B(n82), .Y(n32) );
  INVx1_ASAP7_6t_L U141 ( .A(n83), .Y(n81) );
  INVx1_ASAP7_6t_L U142 ( .A(n80), .Y(n79) );
  XOR2xp5r_ASAP7_6t_L U143 ( .A(n75), .B(n74), .Y(n80) );
  XOR2xp5r_ASAP7_6t_L U144 ( .A(n77), .B(n76), .Y(n74) );
  OAI22xp5_ASAP7_6t_L U145 ( .A1(n84), .A2(n85), .B1(n86), .B2(n87), .Y(n76)
         );
  INVx1_ASAP7_6t_L U146 ( .A(n88), .Y(n84) );
  AO22x1_ASAP7_6t_L U147 ( .A1(n89), .A2(n90), .B1(n59), .B2(n58), .Y(n77) );
  NOR2xp5_ASAP7_6t_L U148 ( .A(n43), .B(n23), .Y(n58) );
  XOR2xp5r_ASAP7_6t_L U149 ( .A(n90), .B(n89), .Y(n59) );
  NOR2xp5_ASAP7_6t_L U150 ( .A(n91), .B(n92), .Y(n90) );
  NOR2xp5_ASAP7_6t_L U151 ( .A(n51), .B(n93), .Y(n89) );
  XOR2xp5r_ASAP7_6t_L U152 ( .A(n94), .B(n95), .Y(n75) );
  OA22x1_ASAP7_6t_L U153 ( .A1(n96), .A2(n97), .B1(n61), .B2(n98), .Y(n78) );
  INVx1_ASAP7_6t_L U154 ( .A(n60), .Y(n98) );
  XOR2xp5r_ASAP7_6t_L U155 ( .A(n97), .B(n96), .Y(n60) );
  XOR2xp5r_ASAP7_6t_L U156 ( .A(n99), .B(n87), .Y(n61) );
  XOR2xp5r_ASAP7_6t_L U157 ( .A(n85), .B(n88), .Y(n87) );
  XOR2xp5r_ASAP7_6t_L U158 ( .A(n100), .B(n101), .Y(n88) );
  INVx1_ASAP7_6t_L U159 ( .A(n102), .Y(n85) );
  NOR3x1f_ASAP7_6t_L U160 ( .A(n103), .B(n24), .C(n49), .Y(n102) );
  INVx1_ASAP7_6t_L U161 ( .A(n86), .Y(n99) );
  XOR2xp5r_ASAP7_6t_L U162 ( .A(n104), .B(n105), .Y(n86) );
  NOR2xp5_ASAP7_6t_L U163 ( .A(n42), .B(n106), .Y(n104) );
  AOI22xp25_ASAP7_6t_L U164 ( .A1(n107), .A2(n108), .B1(n109), .B2(n110), .Y(
        n97) );
  AOI22xp25_ASAP7_6t_L U165 ( .A1(n111), .A2(n112), .B1(n113), .B2(n114), .Y(
        n96) );
  OAI22xp5_ASAP7_6t_L U166 ( .A1(n115), .A2(n116), .B1(n28), .B2(n29), .Y(n242) );
  XOR2xp5r_ASAP7_6t_L U167 ( .A(n116), .B(n117), .Y(n29) );
  XOR2xp5r_ASAP7_6t_L U168 ( .A(n118), .B(n119), .Y(n28) );
  INVx1_ASAP7_6t_L U169 ( .A(n120), .Y(n118) );
  XOR2xp5r_ASAP7_6t_L U170 ( .A(n121), .B(n122), .Y(n116) );
  INVx1_ASAP7_6t_L U171 ( .A(n117), .Y(n115) );
  OAI22xp5_ASAP7_6t_L U172 ( .A1(n123), .A2(n124), .B1(n125), .B2(n72), .Y(
        n117) );
  INVx1_ASAP7_6t_L U173 ( .A(n126), .Y(n72) );
  XOR2xp5r_ASAP7_6t_L U174 ( .A(n127), .B(n128), .Y(n126) );
  INVx1_ASAP7_6t_L U175 ( .A(n73), .Y(n125) );
  XOR2xp5r_ASAP7_6t_L U176 ( .A(n124), .B(n123), .Y(n73) );
  AOI22xp25_ASAP7_6t_L U177 ( .A1(n129), .A2(n130), .B1(n82), .B2(n83), .Y(
        n124) );
  NOR2xp5_ASAP7_6t_L U178 ( .A(n51), .B(n23), .Y(n83) );
  XOR2xp5r_ASAP7_6t_L U179 ( .A(n129), .B(n130), .Y(n82) );
  NOR2xp5_ASAP7_6t_L U180 ( .A(n91), .B(n93), .Y(n130) );
  XOR2xp5r_ASAP7_6t_L U181 ( .A(n131), .B(n132), .Y(n129) );
  NAND2xp5R_ASAP7_6t_L U182 ( .A(a[5]), .B(b[3]), .Y(n131) );
  AOI22xp25_ASAP7_6t_L U183 ( .A1(n133), .A2(n134), .B1(n95), .B2(n94), .Y(
        n123) );
  XOR2xp5r_ASAP7_6t_L U184 ( .A(n133), .B(n134), .Y(n94) );
  XOR2xp5r_ASAP7_6t_L U185 ( .A(n135), .B(n136), .Y(n95) );
  NOR3x1f_ASAP7_6t_L U186 ( .A(n105), .B(n42), .C(n106), .Y(n134) );
  NAND2xp5R_ASAP7_6t_L U187 ( .A(a[3]), .B(b[4]), .Y(n105) );
  AO22x1_ASAP7_6t_L U188 ( .A1(n137), .A2(n138), .B1(n100), .B2(n101), .Y(n133) );
  NOR2xp5_ASAP7_6t_L U189 ( .A(n53), .B(n24), .Y(n101) );
  XOR2xp5r_ASAP7_6t_L U190 ( .A(n138), .B(n137), .Y(n100) );
  NOR2xp5_ASAP7_6t_L U191 ( .A(n52), .B(n50), .Y(n138) );
  NOR2xp5_ASAP7_6t_L U192 ( .A(n49), .B(n139), .Y(n137) );
  AO21x1_ASAP7_6t_L U193 ( .A1(n140), .A2(n141), .B(n142), .Y(n243) );
  NOR3x1f_ASAP7_6t_L U194 ( .A(n143), .B(n23), .C(n27), .Y(n142) );
  INVx1_ASAP7_6t_L U195 ( .A(n26), .Y(n143) );
  XOR2xp5r_ASAP7_6t_L U196 ( .A(n140), .B(n141), .Y(n26) );
  OAI22xp5_ASAP7_6t_L U197 ( .A1(n144), .A2(n145), .B1(n146), .B2(n121), .Y(
        n141) );
  XOR2xp5r_ASAP7_6t_L U198 ( .A(n147), .B(n148), .Y(n121) );
  INVx1_ASAP7_6t_L U199 ( .A(n122), .Y(n146) );
  XOR2xp5r_ASAP7_6t_L U200 ( .A(n145), .B(n144), .Y(n122) );
  AOI22xp25_ASAP7_6t_L U201 ( .A1(n149), .A2(n150), .B1(n71), .B2(n70), .Y(
        n145) );
  NOR2xp5_ASAP7_6t_L U202 ( .A(n91), .B(n23), .Y(n70) );
  XOR2xp5r_ASAP7_6t_L U203 ( .A(n150), .B(n149), .Y(n71) );
  NOR2xp5_ASAP7_6t_L U204 ( .A(n27), .B(n92), .Y(n150) );
  NOR2xp5_ASAP7_6t_L U205 ( .A(n106), .B(n93), .Y(n149) );
  AOI22xp25_ASAP7_6t_L U206 ( .A1(n151), .A2(n152), .B1(n128), .B2(n127), .Y(
        n144) );
  XOR2xp5r_ASAP7_6t_L U207 ( .A(n151), .B(n152), .Y(n127) );
  XOR2xp5r_ASAP7_6t_L U208 ( .A(n153), .B(n154), .Y(n128) );
  NOR3x1f_ASAP7_6t_L U209 ( .A(n132), .B(n92), .C(n106), .Y(n152) );
  NAND2xp5R_ASAP7_6t_L U210 ( .A(b[4]), .B(a[4]), .Y(n132) );
  AO22x1_ASAP7_6t_L U211 ( .A1(n155), .A2(n156), .B1(n135), .B2(n136), .Y(n151) );
  NOR2xp5_ASAP7_6t_L U212 ( .A(n46), .B(n24), .Y(n136) );
  XOR2xp5r_ASAP7_6t_L U213 ( .A(n155), .B(n156), .Y(n135) );
  NOR2xp5_ASAP7_6t_L U214 ( .A(n49), .B(n50), .Y(n156) );
  NOR2xp5_ASAP7_6t_L U215 ( .A(n53), .B(n139), .Y(n155) );
  XOR2xp5r_ASAP7_6t_L U216 ( .A(n157), .B(n158), .Y(n140) );
  AO21x1_ASAP7_6t_L U217 ( .A1(n159), .A2(n160), .B(n161), .Y(n244) );
  NOR3x1f_ASAP7_6t_L U218 ( .A(n24), .B(n162), .C(n23), .Y(n161) );
  INVx1_ASAP7_6t_L U219 ( .A(n22), .Y(n162) );
  XOR2xp5r_ASAP7_6t_L U220 ( .A(n159), .B(n160), .Y(n22) );
  OAI22xp5_ASAP7_6t_L U221 ( .A1(n163), .A2(n164), .B1(n157), .B2(n158), .Y(
        n160) );
  XOR2xp5r_ASAP7_6t_L U222 ( .A(n164), .B(n165), .Y(n158) );
  XOR2xp5r_ASAP7_6t_L U223 ( .A(n166), .B(n167), .Y(n157) );
  INVx1_ASAP7_6t_L U224 ( .A(n168), .Y(n166) );
  AOI22xp25_ASAP7_6t_L U225 ( .A1(n169), .A2(n170), .B1(n120), .B2(n119), .Y(
        n164) );
  NOR2xp5_ASAP7_6t_L U226 ( .A(n106), .B(n23), .Y(n119) );
  XOR2xp5r_ASAP7_6t_L U227 ( .A(n169), .B(n170), .Y(n120) );
  NOR2xp5_ASAP7_6t_L U228 ( .A(n24), .B(n92), .Y(n170) );
  NOR2xp5_ASAP7_6t_L U229 ( .A(n27), .B(n93), .Y(n169) );
  INVx1_ASAP7_6t_L U230 ( .A(n165), .Y(n163) );
  OAI22xp5_ASAP7_6t_L U231 ( .A1(n171), .A2(n172), .B1(n173), .B2(n148), .Y(
        n165) );
  NAND2xp5R_ASAP7_6t_L U232 ( .A(a[4]), .B(b[6]), .Y(n148) );
  INVx1_ASAP7_6t_L U233 ( .A(n147), .Y(n173) );
  XOR2xp5r_ASAP7_6t_L U234 ( .A(n171), .B(n172), .Y(n147) );
  NAND2xp5R_ASAP7_6t_L U235 ( .A(a[3]), .B(b[7]), .Y(n172) );
  AOI22xp25_ASAP7_6t_L U236 ( .A1(n174), .A2(n175), .B1(n153), .B2(n154), .Y(
        n171) );
  NOR2xp5_ASAP7_6t_L U237 ( .A(n42), .B(n24), .Y(n154) );
  XOR2xp5r_ASAP7_6t_L U238 ( .A(n174), .B(n175), .Y(n153) );
  NOR2xp5_ASAP7_6t_L U239 ( .A(n53), .B(n50), .Y(n175) );
  NOR2xp5_ASAP7_6t_L U240 ( .A(n46), .B(n139), .Y(n174) );
  XOR2xp5r_ASAP7_6t_L U241 ( .A(n176), .B(n177), .Y(n159) );
  OR2x2_ASAP7_6t_L U242 ( .A(n178), .B(n179), .Y(n245) );
  NOR3x1f_ASAP7_6t_L U243 ( .A(n50), .B(n180), .C(n93), .Y(n179) );
  NOR3x1f_ASAP7_6t_L U244 ( .A(n20), .B(n23), .C(n139), .Y(n178) );
  INVx1_ASAP7_6t_L U245 ( .A(a[7]), .Y(n23) );
  XOR2xp5r_ASAP7_6t_L U246 ( .A(n181), .B(n180), .Y(n20) );
  OA22x1_ASAP7_6t_L U247 ( .A1(n182), .A2(n183), .B1(n176), .B2(n177), .Y(n180) );
  NAND2xp5R_ASAP7_6t_L U248 ( .A(a[6]), .B(b[6]), .Y(n177) );
  INVx1_ASAP7_6t_L U249 ( .A(n184), .Y(n176) );
  XOR2xp5r_ASAP7_6t_L U250 ( .A(n182), .B(n183), .Y(n184) );
  NAND2xp5R_ASAP7_6t_L U251 ( .A(b[7]), .B(a[5]), .Y(n183) );
  AOI22xp25_ASAP7_6t_L U252 ( .A1(n185), .A2(n186), .B1(n168), .B2(n167), .Y(
        n182) );
  NOR2xp5_ASAP7_6t_L U253 ( .A(n24), .B(n93), .Y(n167) );
  XOR2xp5r_ASAP7_6t_L U254 ( .A(n185), .B(n186), .Y(n168) );
  NOR2xp5_ASAP7_6t_L U255 ( .A(n42), .B(n50), .Y(n186) );
  NOR2xp5_ASAP7_6t_L U256 ( .A(n92), .B(n139), .Y(n185) );
  INVx1_ASAP7_6t_L U257 ( .A(b[6]), .Y(n139) );
  NOR2xp5_ASAP7_6t_L U258 ( .A(n93), .B(n50), .Y(n181) );
  INVx1_ASAP7_6t_L U259 ( .A(b[7]), .Y(n50) );
  INVx1_ASAP7_6t_L U260 ( .A(n273), .Y(n246) );
  INVx1_ASAP7_6t_L U261 ( .A(n272), .Y(out[6]) );
  OAI22xp5_ASAP7_6t_L U262 ( .A1(n187), .A2(n188), .B1(n36), .B2(n37), .Y(n248) );
  XOR2xp5r_ASAP7_6t_L U263 ( .A(n187), .B(n189), .Y(n37) );
  XOR2xp5r_ASAP7_6t_L U264 ( .A(n190), .B(n108), .Y(n36) );
  NOR2xp5_ASAP7_6t_L U265 ( .A(n43), .B(n93), .Y(n108) );
  INVx1_ASAP7_6t_L U266 ( .A(a[6]), .Y(n93) );
  INVx1_ASAP7_6t_L U267 ( .A(n107), .Y(n190) );
  XOR2xp5r_ASAP7_6t_L U268 ( .A(n109), .B(n110), .Y(n107) );
  NOR2xp5_ASAP7_6t_L U269 ( .A(n51), .B(n92), .Y(n110) );
  NOR2xp5_ASAP7_6t_L U270 ( .A(n91), .B(n42), .Y(n109) );
  INVx1_ASAP7_6t_L U271 ( .A(n189), .Y(n188) );
  XOR2xp5r_ASAP7_6t_L U272 ( .A(n63), .B(n62), .Y(n189) );
  XOR2xp5r_ASAP7_6t_L U273 ( .A(n112), .B(n111), .Y(n62) );
  XOR2xp5r_ASAP7_6t_L U274 ( .A(n113), .B(n114), .Y(n111) );
  NOR2xp5_ASAP7_6t_L U275 ( .A(n53), .B(n27), .Y(n114) );
  XOR2xp5r_ASAP7_6t_L U276 ( .A(n103), .B(n191), .Y(n113) );
  NAND2xp5R_ASAP7_6t_L U277 ( .A(a[1]), .B(b[5]), .Y(n191) );
  NAND2xp5R_ASAP7_6t_L U278 ( .A(a[0]), .B(b[6]), .Y(n103) );
  NOR2xp5_ASAP7_6t_L U279 ( .A(n46), .B(n106), .Y(n112) );
  XOR2xp5r_ASAP7_6t_L U280 ( .A(n64), .B(n65), .Y(n63) );
  NOR3x1f_ASAP7_6t_L U281 ( .A(n192), .B(n42), .C(n51), .Y(n65) );
  AO22x1_ASAP7_6t_L U282 ( .A1(n193), .A2(n194), .B1(n195), .B2(n196), .Y(n64)
         );
  AOI22xp25_ASAP7_6t_L U283 ( .A1(n197), .A2(n198), .B1(n199), .B2(n200), .Y(
        n187) );
  INVx1_ASAP7_6t_L U284 ( .A(n271), .Y(n249) );
  INVx1_ASAP7_6t_L U285 ( .A(n270), .Y(out[5]) );
  AO21x1_ASAP7_6t_L U286 ( .A1(n201), .A2(n202), .B(n203), .Y(n251) );
  NOR3x1f_ASAP7_6t_L U287 ( .A(n39), .B(n92), .C(n43), .Y(n203) );
  INVx1_ASAP7_6t_L U288 ( .A(a[5]), .Y(n92) );
  XOR2xp5r_ASAP7_6t_L U289 ( .A(n204), .B(n201), .Y(n39) );
  INVx1_ASAP7_6t_L U290 ( .A(n204), .Y(n202) );
  AOI22xp25_ASAP7_6t_L U291 ( .A1(n205), .A2(n206), .B1(n207), .B2(n208), .Y(
        n204) );
  XOR2xp5r_ASAP7_6t_L U292 ( .A(n198), .B(n197), .Y(n201) );
  XOR2xp5r_ASAP7_6t_L U293 ( .A(n200), .B(n199), .Y(n197) );
  XOR2xp5r_ASAP7_6t_L U294 ( .A(n193), .B(n194), .Y(n199) );
  NOR2xp5_ASAP7_6t_L U295 ( .A(n53), .B(n106), .Y(n194) );
  XOR2xp5r_ASAP7_6t_L U296 ( .A(n195), .B(n196), .Y(n193) );
  NOR2xp5_ASAP7_6t_L U297 ( .A(n49), .B(n27), .Y(n196) );
  INVx1_ASAP7_6t_L U298 ( .A(b[4]), .Y(n27) );
  NOR2xp5_ASAP7_6t_L U299 ( .A(n52), .B(n24), .Y(n195) );
  INVx1_ASAP7_6t_L U300 ( .A(b[5]), .Y(n24) );
  INVx1_ASAP7_6t_L U301 ( .A(a[0]), .Y(n52) );
  NOR3x1f_ASAP7_6t_L U302 ( .A(n209), .B(n106), .C(n49), .Y(n200) );
  INVx1_ASAP7_6t_L U303 ( .A(b[3]), .Y(n106) );
  XOR2xp5r_ASAP7_6t_L U304 ( .A(n210), .B(n192), .Y(n198) );
  NAND2xp5R_ASAP7_6t_L U305 ( .A(b[2]), .B(a[3]), .Y(n192) );
  NAND2xp5R_ASAP7_6t_L U306 ( .A(a[4]), .B(b[1]), .Y(n210) );
  INVx1_ASAP7_6t_L U307 ( .A(n269), .Y(n252) );
  INVx1_ASAP7_6t_L U308 ( .A(n268), .Y(out[4]) );
  AO21x1_ASAP7_6t_L U309 ( .A1(n211), .A2(n212), .B(n213), .Y(n254) );
  NOR3x1f_ASAP7_6t_L U310 ( .A(n43), .B(n214), .C(n42), .Y(n213) );
  INVx1_ASAP7_6t_L U311 ( .A(a[4]), .Y(n42) );
  INVx1_ASAP7_6t_L U312 ( .A(n41), .Y(n214) );
  XOR2xp5r_ASAP7_6t_L U313 ( .A(n212), .B(n211), .Y(n41) );
  XOR2xp5r_ASAP7_6t_L U314 ( .A(n206), .B(n205), .Y(n212) );
  XOR2xp5r_ASAP7_6t_L U315 ( .A(n207), .B(n208), .Y(n205) );
  NOR2xp5_ASAP7_6t_L U316 ( .A(n91), .B(n53), .Y(n208) );
  XOR2xp5r_ASAP7_6t_L U317 ( .A(n209), .B(n215), .Y(n207) );
  NAND2xp5R_ASAP7_6t_L U318 ( .A(a[1]), .B(b[3]), .Y(n215) );
  NAND2xp5R_ASAP7_6t_L U319 ( .A(a[0]), .B(b[4]), .Y(n209) );
  NOR2xp5_ASAP7_6t_L U320 ( .A(n51), .B(n46), .Y(n206) );
  NOR3x1f_ASAP7_6t_L U321 ( .A(n216), .B(n91), .C(n49), .Y(n211) );
  INVx1_ASAP7_6t_L U322 ( .A(n267), .Y(n255) );
  INVx1_ASAP7_6t_L U323 ( .A(n266), .Y(out[3]) );
  OR2x2_ASAP7_6t_L U324 ( .A(n217), .B(n218), .Y(n257) );
  NOR3x1f_ASAP7_6t_L U325 ( .A(n51), .B(n219), .C(n53), .Y(n218) );
  INVx1_ASAP7_6t_L U326 ( .A(a[2]), .Y(n53) );
  NOR3x1f_ASAP7_6t_L U327 ( .A(n43), .B(n220), .C(n46), .Y(n217) );
  INVx1_ASAP7_6t_L U328 ( .A(a[3]), .Y(n46) );
  INVx1_ASAP7_6t_L U329 ( .A(n45), .Y(n220) );
  XOR2xp5r_ASAP7_6t_L U330 ( .A(n219), .B(n221), .Y(n45) );
  NAND2xp5R_ASAP7_6t_L U331 ( .A(b[1]), .B(a[2]), .Y(n221) );
  XOR2xp5r_ASAP7_6t_L U332 ( .A(n222), .B(n216), .Y(n219) );
  NAND2xp5R_ASAP7_6t_L U333 ( .A(a[0]), .B(b[3]), .Y(n216) );
  NOR2xp5_ASAP7_6t_L U334 ( .A(n91), .B(n49), .Y(n222) );
  INVx1_ASAP7_6t_L U335 ( .A(b[2]), .Y(n91) );
  INVx1_ASAP7_6t_L U336 ( .A(b[0]), .Y(n43) );
  INVx1_ASAP7_6t_L U337 ( .A(n265), .Y(n258) );
  INVx1_ASAP7_6t_L U338 ( .A(n264), .Y(out[2]) );
  INVx1_ASAP7_6t_L U339 ( .A(n263), .Y(n260) );
  INVx1_ASAP7_6t_L U340 ( .A(n262), .Y(out[1]) );
  NOR3x1f_ASAP7_6t_L U341 ( .A(n48), .B(n49), .C(n51), .Y(c_30_) );
  INVx1_ASAP7_6t_L U342 ( .A(b[1]), .Y(n51) );
  INVx1_ASAP7_6t_L U343 ( .A(a[1]), .Y(n49) );
  NAND2xp5R_ASAP7_6t_L U344 ( .A(a[0]), .B(b[2]), .Y(n48) );
endmodule

