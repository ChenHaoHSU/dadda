
module DADDA_8x8_42 ( a, b, out );
  input [7:0] a;
  input [7:0] b;
  output [15:0] out;
  wire   n20, n21, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n243, n245, n247, n249, n251, n253, n255,
         n257, n258, n260, n262, n264, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289;
  wire   [63:1] p;
  wire   [23:12] s;
  wire   [22:13] c;

  FAxp33_ASAP7_6t_L add_78_U1_1 ( .A(s[12]), .B(p[16]), .CI(n20), .CON(n267), 
        .SN(n266) );
  FAxp33_ASAP7_6t_L add_78_U1_3 ( .A(s[14]), .B(c[13]), .CI(n21), .CON(n269), 
        .SN(n268) );
  FAxp33_ASAP7_6t_L add_78_U1_4 ( .A(s[15]), .B(c[14]), .CI(n262), .CON(n271), 
        .SN(n270) );
  FAxp33_ASAP7_6t_L add_78_U1_5 ( .A(s[16]), .B(c[15]), .CI(n260), .CON(n273), 
        .SN(n272) );
  FAxp33_ASAP7_6t_L add_78_U1_6 ( .A(s[17]), .B(c[16]), .CI(n258), .CON(n275), 
        .SN(n274) );
  FAxp33_ASAP7_6t_L add_78_U1_7 ( .A(s[18]), .B(c[17]), .CI(n255), .CON(n277), 
        .SN(n276) );
  FAxp33_ASAP7_6t_L add_78_U1_8 ( .A(s[19]), .B(c[18]), .CI(n253), .CON(n279), 
        .SN(n278) );
  FAxp33_ASAP7_6t_L add_78_U1_9 ( .A(s[20]), .B(c[19]), .CI(n251), .CON(n281), 
        .SN(n280) );
  FAxp33_ASAP7_6t_L add_78_U1_10 ( .A(s[21]), .B(c[20]), .CI(n249), .CON(n283), 
        .SN(n282) );
  FAxp33_ASAP7_6t_L add_78_U1_11 ( .A(s[22]), .B(c[21]), .CI(n247), .CON(n285), 
        .SN(n284) );
  FAxp33_ASAP7_6t_L add_78_U1_12 ( .A(s[23]), .B(c[22]), .CI(n245), .CON(n287), 
        .SN(n286) );
  FAxp33_ASAP7_6t_L add_78_U1_13 ( .A(p[63]), .B(n257), .CI(n243), .CON(n289), 
        .SN(n288) );
  AND2x2_ASAP7_6t_L U85 ( .A(p[8]), .B(p[1]), .Y(n20) );
  AND2x2_ASAP7_6t_L U86 ( .A(s[13]), .B(n264), .Y(n21) );
  XOR2xp5r_ASAP7_6t_L U87 ( .A(p[1]), .B(p[8]), .Y(out[1]) );
  XOR2xp5r_ASAP7_6t_L U88 ( .A(n264), .B(s[13]), .Y(out[3]) );
  XOR2xp5r_ASAP7_6t_L U89 ( .A(n24), .B(n25), .Y(s[23]) );
  XOR2xp5r_ASAP7_6t_L U90 ( .A(n26), .B(n27), .Y(s[22]) );
  XOR2xp5r_ASAP7_6t_L U91 ( .A(n28), .B(n29), .Y(s[21]) );
  XOR2xp5r_ASAP7_6t_L U92 ( .A(n30), .B(n31), .Y(s[20]) );
  XOR2xp5r_ASAP7_6t_L U93 ( .A(n32), .B(n33), .Y(s[19]) );
  XOR2xp5r_ASAP7_6t_L U94 ( .A(n34), .B(n35), .Y(s[18]) );
  XOR2xp5r_ASAP7_6t_L U95 ( .A(n36), .B(n37), .Y(s[17]) );
  XOR2xp5r_ASAP7_6t_L U96 ( .A(n38), .B(n39), .Y(s[16]) );
  XOR2xp5r_ASAP7_6t_L U97 ( .A(n40), .B(n41), .Y(s[15]) );
  XOR2xp5r_ASAP7_6t_L U98 ( .A(n42), .B(n43), .Y(s[14]) );
  XOR2xp5r_ASAP7_6t_L U99 ( .A(n44), .B(n45), .Y(s[13]) );
  XOR2xp5r_ASAP7_6t_L U100 ( .A(n46), .B(n47), .Y(s[12]) );
  NAND2xp5R_ASAP7_6t_L U101 ( .A(b[1]), .B(a[1]), .Y(n46) );
  NOR2xp5_ASAP7_6t_L U102 ( .A(n48), .B(n49), .Y(p[8]) );
  NOR2xp5_ASAP7_6t_L U103 ( .A(n50), .B(n51), .Y(p[63]) );
  NOR2xp5_ASAP7_6t_L U104 ( .A(n52), .B(n53), .Y(p[1]) );
  NOR2xp5_ASAP7_6t_L U105 ( .A(n54), .B(n49), .Y(p[16]) );
  NOR2xp5_ASAP7_6t_L U106 ( .A(n52), .B(n49), .Y(out[0]) );
  INVx1_ASAP7_6t_L U107 ( .A(n289), .Y(out[15]) );
  INVx1_ASAP7_6t_L U108 ( .A(n288), .Y(out[14]) );
  INVx1_ASAP7_6t_L U109 ( .A(n287), .Y(n243) );
  INVx1_ASAP7_6t_L U110 ( .A(n286), .Y(out[13]) );
  INVx1_ASAP7_6t_L U111 ( .A(n285), .Y(n245) );
  INVx1_ASAP7_6t_L U112 ( .A(n284), .Y(out[12]) );
  INVx1_ASAP7_6t_L U113 ( .A(n283), .Y(n247) );
  INVx1_ASAP7_6t_L U114 ( .A(n282), .Y(out[11]) );
  INVx1_ASAP7_6t_L U115 ( .A(n281), .Y(n249) );
  INVx1_ASAP7_6t_L U116 ( .A(n280), .Y(out[10]) );
  INVx1_ASAP7_6t_L U117 ( .A(n279), .Y(n251) );
  INVx1_ASAP7_6t_L U118 ( .A(n278), .Y(out[9]) );
  INVx1_ASAP7_6t_L U119 ( .A(n277), .Y(n253) );
  INVx1_ASAP7_6t_L U120 ( .A(n276), .Y(out[8]) );
  INVx1_ASAP7_6t_L U121 ( .A(n275), .Y(n255) );
  INVx1_ASAP7_6t_L U122 ( .A(n274), .Y(out[7]) );
  AO21x1_ASAP7_6t_L U123 ( .A1(n25), .A2(n24), .B(n55), .Y(n257) );
  NOR3x1f_ASAP7_6t_L U124 ( .A(n56), .B(n57), .C(n51), .Y(n55) );
  OR2x2_ASAP7_6t_L U125 ( .A(n58), .B(n59), .Y(n24) );
  NOR3x1f_ASAP7_6t_L U126 ( .A(n60), .B(n61), .C(n50), .Y(n59) );
  NOR3x1f_ASAP7_6t_L U127 ( .A(n62), .B(n57), .C(n63), .Y(n58) );
  XOR2xp5r_ASAP7_6t_L U128 ( .A(n64), .B(n56), .Y(n25) );
  NAND2xp5R_ASAP7_6t_L U129 ( .A(a[6]), .B(b[7]), .Y(n56) );
  NAND2xp5R_ASAP7_6t_L U130 ( .A(b[6]), .B(a[7]), .Y(n64) );
  INVx1_ASAP7_6t_L U131 ( .A(n273), .Y(n258) );
  INVx1_ASAP7_6t_L U132 ( .A(n272), .Y(out[6]) );
  INVx1_ASAP7_6t_L U133 ( .A(n271), .Y(n260) );
  INVx1_ASAP7_6t_L U134 ( .A(n270), .Y(out[5]) );
  INVx1_ASAP7_6t_L U135 ( .A(n269), .Y(n262) );
  INVx1_ASAP7_6t_L U136 ( .A(n268), .Y(out[4]) );
  INVx1_ASAP7_6t_L U137 ( .A(n267), .Y(n264) );
  INVx1_ASAP7_6t_L U138 ( .A(n266), .Y(out[2]) );
  OAI22xp5_ASAP7_6t_L U139 ( .A1(n65), .A2(n66), .B1(n26), .B2(n27), .Y(c[22])
         );
  AOI21xp25_ASAP7_6t_L U140 ( .A1(n67), .A2(n68), .B(n69), .Y(n27) );
  NOR3x1f_ASAP7_6t_L U141 ( .A(n68), .B(n70), .C(n63), .Y(n69) );
  INVx1_ASAP7_6t_L U142 ( .A(n26), .Y(n65) );
  XOR2xp5r_ASAP7_6t_L U143 ( .A(n71), .B(n62), .Y(n26) );
  INVx1_ASAP7_6t_L U144 ( .A(n60), .Y(n62) );
  XOR2xp5r_ASAP7_6t_L U145 ( .A(n72), .B(n73), .Y(n60) );
  NAND2xp5R_ASAP7_6t_L U146 ( .A(b[7]), .B(a[5]), .Y(n73) );
  AOI22xp25_ASAP7_6t_L U147 ( .A1(n74), .A2(n75), .B1(n76), .B2(n77), .Y(n72)
         );
  XOR2xp5r_ASAP7_6t_L U148 ( .A(n78), .B(n66), .Y(n71) );
  NAND2xp5R_ASAP7_6t_L U149 ( .A(a[7]), .B(b[5]), .Y(n66) );
  NAND2xp5R_ASAP7_6t_L U150 ( .A(a[6]), .B(b[6]), .Y(n78) );
  OAI22xp5_ASAP7_6t_L U151 ( .A1(n29), .A2(n28), .B1(n79), .B2(n80), .Y(c[21])
         );
  INVx1_ASAP7_6t_L U152 ( .A(n28), .Y(n79) );
  XOR2xp5r_ASAP7_6t_L U153 ( .A(n81), .B(n68), .Y(n28) );
  AOI22xp25_ASAP7_6t_L U154 ( .A1(n82), .A2(n83), .B1(n84), .B2(n85), .Y(n68)
         );
  XOR2xp5r_ASAP7_6t_L U155 ( .A(n86), .B(n67), .Y(n85) );
  XOR2xp5r_ASAP7_6t_L U156 ( .A(n87), .B(n67), .Y(n83) );
  XOR2xp5r_ASAP7_6t_L U157 ( .A(n77), .B(n76), .Y(n67) );
  AO21x1_ASAP7_6t_L U158 ( .A1(n88), .A2(n89), .B(n90), .Y(n76) );
  NOR3x1f_ASAP7_6t_L U159 ( .A(n89), .B(n61), .C(n70), .Y(n90) );
  XOR2xp5r_ASAP7_6t_L U160 ( .A(n75), .B(n74), .Y(n77) );
  NOR2xp5_ASAP7_6t_L U161 ( .A(n57), .B(n61), .Y(n74) );
  NOR2xp5_ASAP7_6t_L U162 ( .A(n50), .B(n91), .Y(n75) );
  XOR2xp5r_ASAP7_6t_L U163 ( .A(n92), .B(n80), .Y(n81) );
  NAND2xp5R_ASAP7_6t_L U164 ( .A(b[4]), .B(a[7]), .Y(n80) );
  NAND2xp5R_ASAP7_6t_L U165 ( .A(a[6]), .B(b[5]), .Y(n92) );
  AOI21xp25_ASAP7_6t_L U166 ( .A1(n93), .A2(n94), .B(n95), .Y(n29) );
  NOR3x1f_ASAP7_6t_L U167 ( .A(n94), .B(n51), .C(n96), .Y(n95) );
  AO22x1_ASAP7_6t_L U168 ( .A1(n97), .A2(n98), .B1(n31), .B2(n30), .Y(c[20])
         );
  OAI22xp5_ASAP7_6t_L U169 ( .A1(n99), .A2(n100), .B1(n101), .B2(n102), .Y(n30) );
  INVx1_ASAP7_6t_L U170 ( .A(n102), .Y(n99) );
  INVx1_ASAP7_6t_L U171 ( .A(n31), .Y(n98) );
  XOR2xp5r_ASAP7_6t_L U172 ( .A(n103), .B(n94), .Y(n31) );
  AOI22xp25_ASAP7_6t_L U173 ( .A1(n104), .A2(n105), .B1(n106), .B2(n107), .Y(
        n94) );
  XOR2xp5r_ASAP7_6t_L U174 ( .A(n108), .B(n93), .Y(n107) );
  XOR2xp5r_ASAP7_6t_L U175 ( .A(n109), .B(n93), .Y(n105) );
  XOR2xp5r_ASAP7_6t_L U176 ( .A(n82), .B(n87), .Y(n93) );
  AO21x1_ASAP7_6t_L U177 ( .A1(n110), .A2(n111), .B(n112), .Y(n87) );
  NOR3x1f_ASAP7_6t_L U178 ( .A(n111), .B(n91), .C(n70), .Y(n112) );
  INVx1_ASAP7_6t_L U179 ( .A(n84), .Y(n82) );
  XOR2xp5r_ASAP7_6t_L U180 ( .A(n89), .B(n113), .Y(n84) );
  XOR2xp5r_ASAP7_6t_L U181 ( .A(n114), .B(n86), .Y(n113) );
  NOR2xp5_ASAP7_6t_L U182 ( .A(n115), .B(n63), .Y(n86) );
  NOR2xp5_ASAP7_6t_L U183 ( .A(n61), .B(n70), .Y(n114) );
  XOR2xp5r_ASAP7_6t_L U184 ( .A(n116), .B(n88), .Y(n89) );
  NOR2xp5_ASAP7_6t_L U185 ( .A(n117), .B(n50), .Y(n88) );
  NAND2xp5R_ASAP7_6t_L U186 ( .A(b[6]), .B(a[4]), .Y(n116) );
  INVx1_ASAP7_6t_L U187 ( .A(n106), .Y(n104) );
  XOR2xp5r_ASAP7_6t_L U188 ( .A(n118), .B(n97), .Y(n103) );
  NAND2xp5R_ASAP7_6t_L U189 ( .A(b[3]), .B(a[7]), .Y(n118) );
  OAI22xp5_ASAP7_6t_L U190 ( .A1(n119), .A2(n120), .B1(n121), .B2(n122), .Y(
        n97) );
  INVx1_ASAP7_6t_L U191 ( .A(n123), .Y(n120) );
  AO21x1_ASAP7_6t_L U192 ( .A1(n32), .A2(n33), .B(n124), .Y(c[19]) );
  NOR3x1f_ASAP7_6t_L U193 ( .A(n33), .B(n125), .C(n126), .Y(n124) );
  XOR2xp5r_ASAP7_6t_L U194 ( .A(n127), .B(n102), .Y(n33) );
  AOI22xp25_ASAP7_6t_L U195 ( .A1(n128), .A2(n129), .B1(n130), .B2(n131), .Y(
        n102) );
  XOR2xp5r_ASAP7_6t_L U196 ( .A(n132), .B(n100), .Y(n131) );
  INVx1_ASAP7_6t_L U197 ( .A(n128), .Y(n130) );
  XOR2xp5r_ASAP7_6t_L U198 ( .A(n133), .B(n100), .Y(n129) );
  XOR2xp5r_ASAP7_6t_L U199 ( .A(n106), .B(n109), .Y(n100) );
  AO21x1_ASAP7_6t_L U200 ( .A1(n134), .A2(n135), .B(n136), .Y(n109) );
  NOR3x1f_ASAP7_6t_L U201 ( .A(n135), .B(n117), .C(n70), .Y(n136) );
  XOR2xp5r_ASAP7_6t_L U202 ( .A(n111), .B(n137), .Y(n106) );
  XOR2xp5r_ASAP7_6t_L U203 ( .A(n138), .B(n108), .Y(n137) );
  NOR2xp5_ASAP7_6t_L U204 ( .A(n115), .B(n61), .Y(n108) );
  NOR2xp5_ASAP7_6t_L U205 ( .A(n91), .B(n70), .Y(n138) );
  XOR2xp5r_ASAP7_6t_L U206 ( .A(n139), .B(n110), .Y(n111) );
  NOR2xp5_ASAP7_6t_L U207 ( .A(n54), .B(n50), .Y(n110) );
  NAND2xp5R_ASAP7_6t_L U208 ( .A(b[6]), .B(a[3]), .Y(n139) );
  XOR2xp5r_ASAP7_6t_L U209 ( .A(n140), .B(n101), .Y(n127) );
  XOR2xp5r_ASAP7_6t_L U210 ( .A(n119), .B(n123), .Y(n101) );
  XOR2xp5r_ASAP7_6t_L U211 ( .A(n121), .B(n122), .Y(n123) );
  NAND2xp5R_ASAP7_6t_L U212 ( .A(b[3]), .B(a[6]), .Y(n122) );
  NAND2xp5R_ASAP7_6t_L U213 ( .A(b[2]), .B(a[7]), .Y(n121) );
  AOI21xp25_ASAP7_6t_L U214 ( .A1(n141), .A2(n142), .B(n143), .Y(n119) );
  NOR2xp5_ASAP7_6t_L U215 ( .A(n125), .B(n126), .Y(n140) );
  INVx1_ASAP7_6t_L U216 ( .A(n144), .Y(n126) );
  OAI22xp5_ASAP7_6t_L U217 ( .A1(n145), .A2(n146), .B1(n147), .B2(n148), .Y(
        n32) );
  OAI22xp5_ASAP7_6t_L U218 ( .A1(n34), .A2(n35), .B1(n149), .B2(n150), .Y(
        c[18]) );
  INVx1_ASAP7_6t_L U219 ( .A(n149), .Y(n35) );
  XOR2xp5r_ASAP7_6t_L U220 ( .A(n150), .B(n151), .Y(n149) );
  XOR2xp5r_ASAP7_6t_L U221 ( .A(n146), .B(n147), .Y(n151) );
  INVx1_ASAP7_6t_L U222 ( .A(n145), .Y(n147) );
  AOI22xp25_ASAP7_6t_L U223 ( .A1(n152), .A2(n153), .B1(n154), .B2(n155), .Y(
        n145) );
  XOR2xp5r_ASAP7_6t_L U224 ( .A(n156), .B(n148), .Y(n155) );
  INVx1_ASAP7_6t_L U225 ( .A(n152), .Y(n154) );
  XOR2xp5r_ASAP7_6t_L U226 ( .A(n157), .B(n148), .Y(n153) );
  XOR2xp5r_ASAP7_6t_L U227 ( .A(n128), .B(n133), .Y(n148) );
  AOI21xp25_ASAP7_6t_L U228 ( .A1(n158), .A2(n159), .B(n160), .Y(n133) );
  NOR3x1f_ASAP7_6t_L U229 ( .A(n159), .B(n70), .C(n54), .Y(n160) );
  XOR2xp5r_ASAP7_6t_L U230 ( .A(n135), .B(n161), .Y(n128) );
  XOR2xp5r_ASAP7_6t_L U231 ( .A(n162), .B(n132), .Y(n161) );
  NAND2xp5R_ASAP7_6t_L U232 ( .A(b[4]), .B(a[4]), .Y(n132) );
  NOR2xp5_ASAP7_6t_L U233 ( .A(n117), .B(n70), .Y(n162) );
  XOR2xp5r_ASAP7_6t_L U234 ( .A(n163), .B(n134), .Y(n135) );
  NOR2xp5_ASAP7_6t_L U235 ( .A(n48), .B(n50), .Y(n134) );
  NAND2xp5R_ASAP7_6t_L U236 ( .A(b[6]), .B(a[2]), .Y(n163) );
  XOR2xp5r_ASAP7_6t_L U237 ( .A(n144), .B(n125), .Y(n146) );
  AOI21xp25_ASAP7_6t_L U238 ( .A1(n164), .A2(n165), .B(n166), .Y(n125) );
  NOR3x1f_ASAP7_6t_L U239 ( .A(n165), .B(n63), .C(n53), .Y(n166) );
  O2A1O1Ixp33_ASAP7_6t_L U240 ( .A1(n53), .A2(n51), .B(n142), .C(n143), .Y(
        n144) );
  NOR3x1f_ASAP7_6t_L U241 ( .A(n53), .B(n142), .C(n51), .Y(n143) );
  XOR2xp5r_ASAP7_6t_L U242 ( .A(n167), .B(n141), .Y(n142) );
  NOR2xp5_ASAP7_6t_L U243 ( .A(n96), .B(n61), .Y(n141) );
  NAND2xp5R_ASAP7_6t_L U244 ( .A(a[6]), .B(b[2]), .Y(n167) );
  AOI22xp25_ASAP7_6t_L U245 ( .A1(n168), .A2(n169), .B1(n170), .B2(n171), .Y(
        n150) );
  AOI22xp25_ASAP7_6t_L U246 ( .A1(n172), .A2(n173), .B1(n174), .B2(n175), .Y(
        n34) );
  INVx1_ASAP7_6t_L U247 ( .A(n176), .Y(n175) );
  NOR2xp5_ASAP7_6t_L U248 ( .A(n36), .B(n37), .Y(c[17]) );
  XOR2xp5r_ASAP7_6t_L U249 ( .A(n173), .B(n174), .Y(n37) );
  INVx1_ASAP7_6t_L U250 ( .A(n172), .Y(n174) );
  OAI22xp5_ASAP7_6t_L U251 ( .A1(n177), .A2(n178), .B1(n179), .B2(n180), .Y(
        n172) );
  XOR2xp5r_ASAP7_6t_L U252 ( .A(n181), .B(n176), .Y(n180) );
  INVx1_ASAP7_6t_L U253 ( .A(n177), .Y(n179) );
  XOR2xp5r_ASAP7_6t_L U254 ( .A(n182), .B(n176), .Y(n178) );
  XOR2xp5r_ASAP7_6t_L U255 ( .A(n152), .B(n157), .Y(n176) );
  AOI21xp25_ASAP7_6t_L U256 ( .A1(n183), .A2(n184), .B(n185), .Y(n157) );
  NOR3x1f_ASAP7_6t_L U257 ( .A(n184), .B(n54), .C(n115), .Y(n185) );
  XOR2xp5r_ASAP7_6t_L U258 ( .A(n159), .B(n186), .Y(n152) );
  XOR2xp5r_ASAP7_6t_L U259 ( .A(n187), .B(n156), .Y(n186) );
  NAND2xp5R_ASAP7_6t_L U260 ( .A(b[4]), .B(a[3]), .Y(n156) );
  NOR2xp5_ASAP7_6t_L U261 ( .A(n70), .B(n54), .Y(n187) );
  XOR2xp5r_ASAP7_6t_L U262 ( .A(n188), .B(n158), .Y(n159) );
  NOR2xp5_ASAP7_6t_L U263 ( .A(n52), .B(n50), .Y(n158) );
  INVx1_ASAP7_6t_L U264 ( .A(b[7]), .Y(n50) );
  NAND2xp5R_ASAP7_6t_L U265 ( .A(b[6]), .B(a[1]), .Y(n188) );
  XOR2xp5r_ASAP7_6t_L U266 ( .A(n168), .B(n169), .Y(n173) );
  NOR3x1f_ASAP7_6t_L U267 ( .A(n189), .B(n61), .C(n53), .Y(n169) );
  INVx1_ASAP7_6t_L U268 ( .A(n170), .Y(n168) );
  XOR2xp5r_ASAP7_6t_L U269 ( .A(n165), .B(n190), .Y(n170) );
  XOR2xp5r_ASAP7_6t_L U270 ( .A(n191), .B(n171), .Y(n190) );
  NOR2xp5_ASAP7_6t_L U271 ( .A(n49), .B(n51), .Y(n171) );
  INVx1_ASAP7_6t_L U272 ( .A(a[7]), .Y(n51) );
  NOR2xp5_ASAP7_6t_L U273 ( .A(n63), .B(n53), .Y(n191) );
  XOR2xp5r_ASAP7_6t_L U274 ( .A(n192), .B(n164), .Y(n165) );
  NOR2xp5_ASAP7_6t_L U275 ( .A(n96), .B(n91), .Y(n164) );
  INVx1_ASAP7_6t_L U276 ( .A(a[4]), .Y(n91) );
  NAND2xp5R_ASAP7_6t_L U277 ( .A(a[5]), .B(b[2]), .Y(n192) );
  AOI22xp25_ASAP7_6t_L U278 ( .A1(n193), .A2(n194), .B1(n195), .B2(n196), .Y(
        n36) );
  INVx1_ASAP7_6t_L U279 ( .A(n197), .Y(n196) );
  INVx1_ASAP7_6t_L U280 ( .A(n193), .Y(n195) );
  AO21x1_ASAP7_6t_L U281 ( .A1(n39), .A2(n38), .B(n198), .Y(c[16]) );
  NOR3x1f_ASAP7_6t_L U282 ( .A(n39), .B(n63), .C(n49), .Y(n198) );
  AO21x1_ASAP7_6t_L U283 ( .A1(n199), .A2(n200), .B(n201), .Y(n38) );
  XOR2xp5r_ASAP7_6t_L U284 ( .A(n202), .B(n193), .Y(n39) );
  OAI22xp5_ASAP7_6t_L U285 ( .A1(n203), .A2(n204), .B1(n205), .B2(n206), .Y(
        n193) );
  XOR2xp5r_ASAP7_6t_L U286 ( .A(n207), .B(n197), .Y(n206) );
  XOR2xp5r_ASAP7_6t_L U287 ( .A(n208), .B(n197), .Y(n204) );
  XOR2xp5r_ASAP7_6t_L U288 ( .A(n177), .B(n182), .Y(n197) );
  AO21x1_ASAP7_6t_L U289 ( .A1(n209), .A2(n210), .B(n211), .Y(n182) );
  NOR3x1f_ASAP7_6t_L U290 ( .A(n210), .B(n54), .C(n96), .Y(n211) );
  XOR2xp5r_ASAP7_6t_L U291 ( .A(n184), .B(n212), .Y(n177) );
  XOR2xp5r_ASAP7_6t_L U292 ( .A(n213), .B(n181), .Y(n212) );
  NOR2xp5_ASAP7_6t_L U293 ( .A(n96), .B(n117), .Y(n181) );
  NOR2xp5_ASAP7_6t_L U294 ( .A(n54), .B(n115), .Y(n213) );
  INVx1_ASAP7_6t_L U295 ( .A(b[4]), .Y(n115) );
  XOR2xp5r_ASAP7_6t_L U296 ( .A(n214), .B(n183), .Y(n184) );
  NOR2xp5_ASAP7_6t_L U297 ( .A(n52), .B(n57), .Y(n183) );
  INVx1_ASAP7_6t_L U298 ( .A(b[6]), .Y(n57) );
  NAND2xp5R_ASAP7_6t_L U299 ( .A(b[5]), .B(a[1]), .Y(n214) );
  XOR2xp5r_ASAP7_6t_L U300 ( .A(n215), .B(n194), .Y(n202) );
  XOR2xp5r_ASAP7_6t_L U301 ( .A(n189), .B(n216), .Y(n194) );
  NAND2xp5R_ASAP7_6t_L U302 ( .A(b[1]), .B(a[5]), .Y(n216) );
  NAND2xp5R_ASAP7_6t_L U303 ( .A(b[2]), .B(a[4]), .Y(n189) );
  NOR2xp5_ASAP7_6t_L U304 ( .A(n63), .B(n49), .Y(n215) );
  INVx1_ASAP7_6t_L U305 ( .A(a[6]), .Y(n63) );
  NOR2xp5_ASAP7_6t_L U306 ( .A(n41), .B(n40), .Y(c[15]) );
  INVx1_ASAP7_6t_L U307 ( .A(n217), .Y(n40) );
  O2A1O1Ixp33_ASAP7_6t_L U308 ( .A1(n49), .A2(n61), .B(n200), .C(n201), .Y(
        n217) );
  NOR3x1f_ASAP7_6t_L U309 ( .A(n49), .B(n200), .C(n61), .Y(n201) );
  XOR2xp5r_ASAP7_6t_L U310 ( .A(n218), .B(n199), .Y(n200) );
  XOR2xp5r_ASAP7_6t_L U311 ( .A(n205), .B(n208), .Y(n199) );
  NOR3x1f_ASAP7_6t_L U312 ( .A(n219), .B(n48), .C(n96), .Y(n208) );
  INVx1_ASAP7_6t_L U313 ( .A(n203), .Y(n205) );
  XOR2xp5r_ASAP7_6t_L U314 ( .A(n210), .B(n220), .Y(n203) );
  XOR2xp5r_ASAP7_6t_L U315 ( .A(n221), .B(n207), .Y(n220) );
  AND2x2_ASAP7_6t_L U316 ( .A(b[2]), .B(a[3]), .Y(n207) );
  NOR2xp5_ASAP7_6t_L U317 ( .A(n54), .B(n96), .Y(n221) );
  XOR2xp5r_ASAP7_6t_L U318 ( .A(n222), .B(n209), .Y(n210) );
  NOR2xp5_ASAP7_6t_L U319 ( .A(n52), .B(n70), .Y(n209) );
  INVx1_ASAP7_6t_L U320 ( .A(b[5]), .Y(n70) );
  NAND2xp5R_ASAP7_6t_L U321 ( .A(b[4]), .B(a[1]), .Y(n222) );
  NAND2xp5R_ASAP7_6t_L U322 ( .A(a[4]), .B(b[1]), .Y(n218) );
  INVx1_ASAP7_6t_L U323 ( .A(a[5]), .Y(n61) );
  INVx1_ASAP7_6t_L U324 ( .A(b[0]), .Y(n49) );
  AOI21xp25_ASAP7_6t_L U325 ( .A1(n223), .A2(n224), .B(n225), .Y(n41) );
  NOR3x1f_ASAP7_6t_L U326 ( .A(n224), .B(n117), .C(n53), .Y(n225) );
  INVx1_ASAP7_6t_L U327 ( .A(a[3]), .Y(n117) );
  OAI22xp5_ASAP7_6t_L U328 ( .A1(n43), .A2(n42), .B1(n226), .B2(n227), .Y(
        c[14]) );
  INVx1_ASAP7_6t_L U329 ( .A(n42), .Y(n226) );
  XOR2xp5r_ASAP7_6t_L U330 ( .A(n228), .B(n224), .Y(n42) );
  XOR2xp5r_ASAP7_6t_L U331 ( .A(n223), .B(n229), .Y(n224) );
  NAND2xp5R_ASAP7_6t_L U332 ( .A(b[2]), .B(a[2]), .Y(n229) );
  XOR2xp5r_ASAP7_6t_L U333 ( .A(n230), .B(n219), .Y(n223) );
  NAND2xp5R_ASAP7_6t_L U334 ( .A(a[0]), .B(b[4]), .Y(n219) );
  NAND2xp5R_ASAP7_6t_L U335 ( .A(a[1]), .B(b[3]), .Y(n230) );
  XOR2xp5r_ASAP7_6t_L U336 ( .A(n231), .B(n227), .Y(n228) );
  NAND2xp5R_ASAP7_6t_L U337 ( .A(b[0]), .B(a[4]), .Y(n227) );
  NAND2xp5R_ASAP7_6t_L U338 ( .A(b[1]), .B(a[3]), .Y(n231) );
  AOI21xp25_ASAP7_6t_L U339 ( .A1(n232), .A2(n233), .B(n234), .Y(n43) );
  NOR3x1f_ASAP7_6t_L U340 ( .A(n233), .B(n54), .C(n53), .Y(n234) );
  INVx1_ASAP7_6t_L U341 ( .A(a[2]), .Y(n54) );
  OAI22xp5_ASAP7_6t_L U342 ( .A1(n45), .A2(n44), .B1(n235), .B2(n236), .Y(
        c[13]) );
  INVx1_ASAP7_6t_L U343 ( .A(n45), .Y(n235) );
  INVx1_ASAP7_6t_L U344 ( .A(n237), .Y(n44) );
  NOR3x1f_ASAP7_6t_L U345 ( .A(n47), .B(n48), .C(n53), .Y(n237) );
  INVx1_ASAP7_6t_L U346 ( .A(b[1]), .Y(n53) );
  INVx1_ASAP7_6t_L U347 ( .A(a[1]), .Y(n48) );
  NAND2xp5R_ASAP7_6t_L U348 ( .A(b[2]), .B(a[0]), .Y(n47) );
  XOR2xp5r_ASAP7_6t_L U349 ( .A(n238), .B(n233), .Y(n45) );
  XOR2xp5r_ASAP7_6t_L U350 ( .A(n239), .B(n232), .Y(n233) );
  NOR2xp5_ASAP7_6t_L U351 ( .A(n52), .B(n96), .Y(n232) );
  INVx1_ASAP7_6t_L U352 ( .A(b[3]), .Y(n96) );
  INVx1_ASAP7_6t_L U353 ( .A(a[0]), .Y(n52) );
  NAND2xp5R_ASAP7_6t_L U354 ( .A(a[1]), .B(b[2]), .Y(n239) );
  XOR2xp5r_ASAP7_6t_L U355 ( .A(n240), .B(n236), .Y(n238) );
  NAND2xp5R_ASAP7_6t_L U356 ( .A(b[0]), .B(a[3]), .Y(n236) );
  NAND2xp5R_ASAP7_6t_L U357 ( .A(b[1]), .B(a[2]), .Y(n240) );
endmodule

